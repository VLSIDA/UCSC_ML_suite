VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_1x256_1r1w
  FOREIGN fakeram_1x256_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 5.184 BY 20.736 ;
  CLASS BLOCK ;
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.276 0.024 0.300 ;
    END
  END w0_wd_in[0]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 0.000 0.225 0.018 ;
    END
  END r0_rd_out[0]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.484 0.024 2.508 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.692 0.024 4.716 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.900 0.024 6.924 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.108 0.024 9.132 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 5.160 0.276 5.184 0.300 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 5.160 2.484 5.184 2.508 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 5.160 4.692 5.184 4.716 ;
    END
  END w0_addr_in[6]
  PIN w0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 5.160 6.900 5.184 6.924 ;
    END
  END w0_addr_in[7]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.316 0.024 11.340 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.524 0.024 13.548 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.732 0.024 15.756 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.940 0.024 17.964 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 5.160 9.108 5.184 9.132 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 5.160 11.316 5.184 11.340 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 5.160 13.524 5.184 13.548 ;
    END
  END r0_addr_in[6]
  PIN r0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 5.160 15.732 5.184 15.756 ;
    END
  END r0_addr_in[7]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 20.718 0.225 20.736 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.963 20.718 0.981 20.736 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.719 20.718 1.737 20.736 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.475 20.718 2.493 20.736 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.231 20.718 3.249 20.736 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.108 0.192 5.076 0.288 ;
      RECT 0.108 0.960 5.076 1.056 ;
      RECT 0.108 1.728 5.076 1.824 ;
      RECT 0.108 2.496 5.076 2.592 ;
      RECT 0.108 3.264 5.076 3.360 ;
      RECT 0.108 4.032 5.076 4.128 ;
      RECT 0.108 4.800 5.076 4.896 ;
      RECT 0.108 5.568 5.076 5.664 ;
      RECT 0.108 6.336 5.076 6.432 ;
      RECT 0.108 7.104 5.076 7.200 ;
      RECT 0.108 7.872 5.076 7.968 ;
      RECT 0.108 8.640 5.076 8.736 ;
      RECT 0.108 9.408 5.076 9.504 ;
      RECT 0.108 10.176 5.076 10.272 ;
      RECT 0.108 10.944 5.076 11.040 ;
      RECT 0.108 11.712 5.076 11.808 ;
      RECT 0.108 12.480 5.076 12.576 ;
      RECT 0.108 13.248 5.076 13.344 ;
      RECT 0.108 14.016 5.076 14.112 ;
      RECT 0.108 14.784 5.076 14.880 ;
      RECT 0.108 15.552 5.076 15.648 ;
      RECT 0.108 16.320 5.076 16.416 ;
      RECT 0.108 17.088 5.076 17.184 ;
      RECT 0.108 17.856 5.076 17.952 ;
      RECT 0.108 18.624 5.076 18.720 ;
      RECT 0.108 19.392 5.076 19.488 ;
      RECT 0.108 20.160 5.076 20.256 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.108 0.192 5.076 0.288 ;
      RECT 0.108 0.960 5.076 1.056 ;
      RECT 0.108 1.728 5.076 1.824 ;
      RECT 0.108 2.496 5.076 2.592 ;
      RECT 0.108 3.264 5.076 3.360 ;
      RECT 0.108 4.032 5.076 4.128 ;
      RECT 0.108 4.800 5.076 4.896 ;
      RECT 0.108 5.568 5.076 5.664 ;
      RECT 0.108 6.336 5.076 6.432 ;
      RECT 0.108 7.104 5.076 7.200 ;
      RECT 0.108 7.872 5.076 7.968 ;
      RECT 0.108 8.640 5.076 8.736 ;
      RECT 0.108 9.408 5.076 9.504 ;
      RECT 0.108 10.176 5.076 10.272 ;
      RECT 0.108 10.944 5.076 11.040 ;
      RECT 0.108 11.712 5.076 11.808 ;
      RECT 0.108 12.480 5.076 12.576 ;
      RECT 0.108 13.248 5.076 13.344 ;
      RECT 0.108 14.016 5.076 14.112 ;
      RECT 0.108 14.784 5.076 14.880 ;
      RECT 0.108 15.552 5.076 15.648 ;
      RECT 0.108 16.320 5.076 16.416 ;
      RECT 0.108 17.088 5.076 17.184 ;
      RECT 0.108 17.856 5.076 17.952 ;
      RECT 0.108 18.624 5.076 18.720 ;
      RECT 0.108 19.392 5.076 19.488 ;
      RECT 0.108 20.160 5.076 20.256 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 5.184 20.736 ;
    LAYER M2 ;
    RECT 0 0 5.184 20.736 ;
    LAYER M3 ;
    RECT 0 0 5.184 20.736 ;
    LAYER M4 ;
    RECT 0 0 5.184 20.736 ;
  END
END fakeram_1x256_1r1w

END LIBRARY
