VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_512x2048_1r1w
  FOREIGN fakeram_512x2048_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 265.421 BY 165.888 ;
  CLASS BLOCK ;
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.276 0.024 0.300 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.428 0.024 1.452 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.580 0.024 2.604 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.732 0.024 3.756 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.884 0.024 4.908 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.036 0.024 6.060 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.188 0.024 7.212 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.340 0.024 8.364 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.492 0.024 9.516 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.644 0.024 10.668 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.796 0.024 11.820 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.948 0.024 12.972 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.100 0.024 14.124 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.252 0.024 15.276 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.404 0.024 16.428 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.556 0.024 17.580 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.708 0.024 18.732 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.860 0.024 19.884 ;
    END
  END w0_wd_in[17]
  PIN w0_wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.012 0.024 21.036 ;
    END
  END w0_wd_in[18]
  PIN w0_wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.164 0.024 22.188 ;
    END
  END w0_wd_in[19]
  PIN w0_wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.316 0.024 23.340 ;
    END
  END w0_wd_in[20]
  PIN w0_wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.468 0.024 24.492 ;
    END
  END w0_wd_in[21]
  PIN w0_wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.620 0.024 25.644 ;
    END
  END w0_wd_in[22]
  PIN w0_wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.772 0.024 26.796 ;
    END
  END w0_wd_in[23]
  PIN w0_wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.924 0.024 27.948 ;
    END
  END w0_wd_in[24]
  PIN w0_wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.076 0.024 29.100 ;
    END
  END w0_wd_in[25]
  PIN w0_wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.228 0.024 30.252 ;
    END
  END w0_wd_in[26]
  PIN w0_wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.380 0.024 31.404 ;
    END
  END w0_wd_in[27]
  PIN w0_wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.532 0.024 32.556 ;
    END
  END w0_wd_in[28]
  PIN w0_wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 33.684 0.024 33.708 ;
    END
  END w0_wd_in[29]
  PIN w0_wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 34.836 0.024 34.860 ;
    END
  END w0_wd_in[30]
  PIN w0_wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 35.988 0.024 36.012 ;
    END
  END w0_wd_in[31]
  PIN w0_wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 37.140 0.024 37.164 ;
    END
  END w0_wd_in[32]
  PIN w0_wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 38.292 0.024 38.316 ;
    END
  END w0_wd_in[33]
  PIN w0_wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 39.444 0.024 39.468 ;
    END
  END w0_wd_in[34]
  PIN w0_wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 40.596 0.024 40.620 ;
    END
  END w0_wd_in[35]
  PIN w0_wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 41.748 0.024 41.772 ;
    END
  END w0_wd_in[36]
  PIN w0_wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 42.900 0.024 42.924 ;
    END
  END w0_wd_in[37]
  PIN w0_wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 44.052 0.024 44.076 ;
    END
  END w0_wd_in[38]
  PIN w0_wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 45.204 0.024 45.228 ;
    END
  END w0_wd_in[39]
  PIN w0_wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 46.356 0.024 46.380 ;
    END
  END w0_wd_in[40]
  PIN w0_wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 47.508 0.024 47.532 ;
    END
  END w0_wd_in[41]
  PIN w0_wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 48.660 0.024 48.684 ;
    END
  END w0_wd_in[42]
  PIN w0_wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 49.812 0.024 49.836 ;
    END
  END w0_wd_in[43]
  PIN w0_wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 50.964 0.024 50.988 ;
    END
  END w0_wd_in[44]
  PIN w0_wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 52.116 0.024 52.140 ;
    END
  END w0_wd_in[45]
  PIN w0_wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 53.268 0.024 53.292 ;
    END
  END w0_wd_in[46]
  PIN w0_wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 54.420 0.024 54.444 ;
    END
  END w0_wd_in[47]
  PIN w0_wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 55.572 0.024 55.596 ;
    END
  END w0_wd_in[48]
  PIN w0_wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 56.724 0.024 56.748 ;
    END
  END w0_wd_in[49]
  PIN w0_wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 57.876 0.024 57.900 ;
    END
  END w0_wd_in[50]
  PIN w0_wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 59.028 0.024 59.052 ;
    END
  END w0_wd_in[51]
  PIN w0_wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 60.180 0.024 60.204 ;
    END
  END w0_wd_in[52]
  PIN w0_wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 61.332 0.024 61.356 ;
    END
  END w0_wd_in[53]
  PIN w0_wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 62.484 0.024 62.508 ;
    END
  END w0_wd_in[54]
  PIN w0_wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 63.636 0.024 63.660 ;
    END
  END w0_wd_in[55]
  PIN w0_wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 64.788 0.024 64.812 ;
    END
  END w0_wd_in[56]
  PIN w0_wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 65.940 0.024 65.964 ;
    END
  END w0_wd_in[57]
  PIN w0_wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 67.092 0.024 67.116 ;
    END
  END w0_wd_in[58]
  PIN w0_wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 68.244 0.024 68.268 ;
    END
  END w0_wd_in[59]
  PIN w0_wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 69.396 0.024 69.420 ;
    END
  END w0_wd_in[60]
  PIN w0_wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 70.548 0.024 70.572 ;
    END
  END w0_wd_in[61]
  PIN w0_wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 71.700 0.024 71.724 ;
    END
  END w0_wd_in[62]
  PIN w0_wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 72.852 0.024 72.876 ;
    END
  END w0_wd_in[63]
  PIN w0_wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 74.004 0.024 74.028 ;
    END
  END w0_wd_in[64]
  PIN w0_wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 75.156 0.024 75.180 ;
    END
  END w0_wd_in[65]
  PIN w0_wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 76.308 0.024 76.332 ;
    END
  END w0_wd_in[66]
  PIN w0_wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 77.460 0.024 77.484 ;
    END
  END w0_wd_in[67]
  PIN w0_wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 78.612 0.024 78.636 ;
    END
  END w0_wd_in[68]
  PIN w0_wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 79.764 0.024 79.788 ;
    END
  END w0_wd_in[69]
  PIN w0_wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 80.916 0.024 80.940 ;
    END
  END w0_wd_in[70]
  PIN w0_wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 82.068 0.024 82.092 ;
    END
  END w0_wd_in[71]
  PIN w0_wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 83.220 0.024 83.244 ;
    END
  END w0_wd_in[72]
  PIN w0_wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 84.372 0.024 84.396 ;
    END
  END w0_wd_in[73]
  PIN w0_wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 85.524 0.024 85.548 ;
    END
  END w0_wd_in[74]
  PIN w0_wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 86.676 0.024 86.700 ;
    END
  END w0_wd_in[75]
  PIN w0_wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 87.828 0.024 87.852 ;
    END
  END w0_wd_in[76]
  PIN w0_wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 88.980 0.024 89.004 ;
    END
  END w0_wd_in[77]
  PIN w0_wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 90.132 0.024 90.156 ;
    END
  END w0_wd_in[78]
  PIN w0_wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 91.284 0.024 91.308 ;
    END
  END w0_wd_in[79]
  PIN w0_wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 92.436 0.024 92.460 ;
    END
  END w0_wd_in[80]
  PIN w0_wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 93.588 0.024 93.612 ;
    END
  END w0_wd_in[81]
  PIN w0_wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 94.740 0.024 94.764 ;
    END
  END w0_wd_in[82]
  PIN w0_wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 95.892 0.024 95.916 ;
    END
  END w0_wd_in[83]
  PIN w0_wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 97.044 0.024 97.068 ;
    END
  END w0_wd_in[84]
  PIN w0_wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 98.196 0.024 98.220 ;
    END
  END w0_wd_in[85]
  PIN w0_wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 99.348 0.024 99.372 ;
    END
  END w0_wd_in[86]
  PIN w0_wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 100.500 0.024 100.524 ;
    END
  END w0_wd_in[87]
  PIN w0_wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 101.652 0.024 101.676 ;
    END
  END w0_wd_in[88]
  PIN w0_wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 102.804 0.024 102.828 ;
    END
  END w0_wd_in[89]
  PIN w0_wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 103.956 0.024 103.980 ;
    END
  END w0_wd_in[90]
  PIN w0_wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 105.108 0.024 105.132 ;
    END
  END w0_wd_in[91]
  PIN w0_wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 106.260 0.024 106.284 ;
    END
  END w0_wd_in[92]
  PIN w0_wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 107.412 0.024 107.436 ;
    END
  END w0_wd_in[93]
  PIN w0_wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 108.564 0.024 108.588 ;
    END
  END w0_wd_in[94]
  PIN w0_wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 109.716 0.024 109.740 ;
    END
  END w0_wd_in[95]
  PIN w0_wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 110.868 0.024 110.892 ;
    END
  END w0_wd_in[96]
  PIN w0_wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 112.020 0.024 112.044 ;
    END
  END w0_wd_in[97]
  PIN w0_wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 113.172 0.024 113.196 ;
    END
  END w0_wd_in[98]
  PIN w0_wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 114.324 0.024 114.348 ;
    END
  END w0_wd_in[99]
  PIN w0_wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 115.476 0.024 115.500 ;
    END
  END w0_wd_in[100]
  PIN w0_wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 116.628 0.024 116.652 ;
    END
  END w0_wd_in[101]
  PIN w0_wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 117.780 0.024 117.804 ;
    END
  END w0_wd_in[102]
  PIN w0_wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 118.932 0.024 118.956 ;
    END
  END w0_wd_in[103]
  PIN w0_wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 120.084 0.024 120.108 ;
    END
  END w0_wd_in[104]
  PIN w0_wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 121.236 0.024 121.260 ;
    END
  END w0_wd_in[105]
  PIN w0_wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 122.388 0.024 122.412 ;
    END
  END w0_wd_in[106]
  PIN w0_wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 123.540 0.024 123.564 ;
    END
  END w0_wd_in[107]
  PIN w0_wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 124.692 0.024 124.716 ;
    END
  END w0_wd_in[108]
  PIN w0_wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 125.844 0.024 125.868 ;
    END
  END w0_wd_in[109]
  PIN w0_wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 126.996 0.024 127.020 ;
    END
  END w0_wd_in[110]
  PIN w0_wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 128.148 0.024 128.172 ;
    END
  END w0_wd_in[111]
  PIN w0_wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 129.300 0.024 129.324 ;
    END
  END w0_wd_in[112]
  PIN w0_wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 130.452 0.024 130.476 ;
    END
  END w0_wd_in[113]
  PIN w0_wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 131.604 0.024 131.628 ;
    END
  END w0_wd_in[114]
  PIN w0_wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 132.756 0.024 132.780 ;
    END
  END w0_wd_in[115]
  PIN w0_wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 133.908 0.024 133.932 ;
    END
  END w0_wd_in[116]
  PIN w0_wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 135.060 0.024 135.084 ;
    END
  END w0_wd_in[117]
  PIN w0_wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 136.212 0.024 136.236 ;
    END
  END w0_wd_in[118]
  PIN w0_wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 137.364 0.024 137.388 ;
    END
  END w0_wd_in[119]
  PIN w0_wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 138.516 0.024 138.540 ;
    END
  END w0_wd_in[120]
  PIN w0_wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 139.668 0.024 139.692 ;
    END
  END w0_wd_in[121]
  PIN w0_wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 140.820 0.024 140.844 ;
    END
  END w0_wd_in[122]
  PIN w0_wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 141.972 0.024 141.996 ;
    END
  END w0_wd_in[123]
  PIN w0_wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 143.124 0.024 143.148 ;
    END
  END w0_wd_in[124]
  PIN w0_wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 144.276 0.024 144.300 ;
    END
  END w0_wd_in[125]
  PIN w0_wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 145.428 0.024 145.452 ;
    END
  END w0_wd_in[126]
  PIN w0_wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 146.580 0.024 146.604 ;
    END
  END w0_wd_in[127]
  PIN w0_wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 0.276 265.421 0.300 ;
    END
  END w0_wd_in[128]
  PIN w0_wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 1.428 265.421 1.452 ;
    END
  END w0_wd_in[129]
  PIN w0_wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 2.580 265.421 2.604 ;
    END
  END w0_wd_in[130]
  PIN w0_wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 3.732 265.421 3.756 ;
    END
  END w0_wd_in[131]
  PIN w0_wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 4.884 265.421 4.908 ;
    END
  END w0_wd_in[132]
  PIN w0_wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 6.036 265.421 6.060 ;
    END
  END w0_wd_in[133]
  PIN w0_wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 7.188 265.421 7.212 ;
    END
  END w0_wd_in[134]
  PIN w0_wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 8.340 265.421 8.364 ;
    END
  END w0_wd_in[135]
  PIN w0_wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 9.492 265.421 9.516 ;
    END
  END w0_wd_in[136]
  PIN w0_wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 10.644 265.421 10.668 ;
    END
  END w0_wd_in[137]
  PIN w0_wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 11.796 265.421 11.820 ;
    END
  END w0_wd_in[138]
  PIN w0_wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 12.948 265.421 12.972 ;
    END
  END w0_wd_in[139]
  PIN w0_wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 14.100 265.421 14.124 ;
    END
  END w0_wd_in[140]
  PIN w0_wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 15.252 265.421 15.276 ;
    END
  END w0_wd_in[141]
  PIN w0_wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 16.404 265.421 16.428 ;
    END
  END w0_wd_in[142]
  PIN w0_wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 17.556 265.421 17.580 ;
    END
  END w0_wd_in[143]
  PIN w0_wd_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 18.708 265.421 18.732 ;
    END
  END w0_wd_in[144]
  PIN w0_wd_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 19.860 265.421 19.884 ;
    END
  END w0_wd_in[145]
  PIN w0_wd_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 21.012 265.421 21.036 ;
    END
  END w0_wd_in[146]
  PIN w0_wd_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 22.164 265.421 22.188 ;
    END
  END w0_wd_in[147]
  PIN w0_wd_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 23.316 265.421 23.340 ;
    END
  END w0_wd_in[148]
  PIN w0_wd_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 24.468 265.421 24.492 ;
    END
  END w0_wd_in[149]
  PIN w0_wd_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 25.620 265.421 25.644 ;
    END
  END w0_wd_in[150]
  PIN w0_wd_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 26.772 265.421 26.796 ;
    END
  END w0_wd_in[151]
  PIN w0_wd_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 27.924 265.421 27.948 ;
    END
  END w0_wd_in[152]
  PIN w0_wd_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 29.076 265.421 29.100 ;
    END
  END w0_wd_in[153]
  PIN w0_wd_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 30.228 265.421 30.252 ;
    END
  END w0_wd_in[154]
  PIN w0_wd_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 31.380 265.421 31.404 ;
    END
  END w0_wd_in[155]
  PIN w0_wd_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 32.532 265.421 32.556 ;
    END
  END w0_wd_in[156]
  PIN w0_wd_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 33.684 265.421 33.708 ;
    END
  END w0_wd_in[157]
  PIN w0_wd_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 34.836 265.421 34.860 ;
    END
  END w0_wd_in[158]
  PIN w0_wd_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 35.988 265.421 36.012 ;
    END
  END w0_wd_in[159]
  PIN w0_wd_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 37.140 265.421 37.164 ;
    END
  END w0_wd_in[160]
  PIN w0_wd_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 38.292 265.421 38.316 ;
    END
  END w0_wd_in[161]
  PIN w0_wd_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 39.444 265.421 39.468 ;
    END
  END w0_wd_in[162]
  PIN w0_wd_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 40.596 265.421 40.620 ;
    END
  END w0_wd_in[163]
  PIN w0_wd_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 41.748 265.421 41.772 ;
    END
  END w0_wd_in[164]
  PIN w0_wd_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 42.900 265.421 42.924 ;
    END
  END w0_wd_in[165]
  PIN w0_wd_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 44.052 265.421 44.076 ;
    END
  END w0_wd_in[166]
  PIN w0_wd_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 45.204 265.421 45.228 ;
    END
  END w0_wd_in[167]
  PIN w0_wd_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 46.356 265.421 46.380 ;
    END
  END w0_wd_in[168]
  PIN w0_wd_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 47.508 265.421 47.532 ;
    END
  END w0_wd_in[169]
  PIN w0_wd_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 48.660 265.421 48.684 ;
    END
  END w0_wd_in[170]
  PIN w0_wd_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 49.812 265.421 49.836 ;
    END
  END w0_wd_in[171]
  PIN w0_wd_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 50.964 265.421 50.988 ;
    END
  END w0_wd_in[172]
  PIN w0_wd_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 52.116 265.421 52.140 ;
    END
  END w0_wd_in[173]
  PIN w0_wd_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 53.268 265.421 53.292 ;
    END
  END w0_wd_in[174]
  PIN w0_wd_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 54.420 265.421 54.444 ;
    END
  END w0_wd_in[175]
  PIN w0_wd_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 55.572 265.421 55.596 ;
    END
  END w0_wd_in[176]
  PIN w0_wd_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 56.724 265.421 56.748 ;
    END
  END w0_wd_in[177]
  PIN w0_wd_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 57.876 265.421 57.900 ;
    END
  END w0_wd_in[178]
  PIN w0_wd_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 59.028 265.421 59.052 ;
    END
  END w0_wd_in[179]
  PIN w0_wd_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 60.180 265.421 60.204 ;
    END
  END w0_wd_in[180]
  PIN w0_wd_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 61.332 265.421 61.356 ;
    END
  END w0_wd_in[181]
  PIN w0_wd_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 62.484 265.421 62.508 ;
    END
  END w0_wd_in[182]
  PIN w0_wd_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 63.636 265.421 63.660 ;
    END
  END w0_wd_in[183]
  PIN w0_wd_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 64.788 265.421 64.812 ;
    END
  END w0_wd_in[184]
  PIN w0_wd_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 65.940 265.421 65.964 ;
    END
  END w0_wd_in[185]
  PIN w0_wd_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 67.092 265.421 67.116 ;
    END
  END w0_wd_in[186]
  PIN w0_wd_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 68.244 265.421 68.268 ;
    END
  END w0_wd_in[187]
  PIN w0_wd_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 69.396 265.421 69.420 ;
    END
  END w0_wd_in[188]
  PIN w0_wd_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 70.548 265.421 70.572 ;
    END
  END w0_wd_in[189]
  PIN w0_wd_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 71.700 265.421 71.724 ;
    END
  END w0_wd_in[190]
  PIN w0_wd_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 72.852 265.421 72.876 ;
    END
  END w0_wd_in[191]
  PIN w0_wd_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 74.004 265.421 74.028 ;
    END
  END w0_wd_in[192]
  PIN w0_wd_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 75.156 265.421 75.180 ;
    END
  END w0_wd_in[193]
  PIN w0_wd_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 76.308 265.421 76.332 ;
    END
  END w0_wd_in[194]
  PIN w0_wd_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 77.460 265.421 77.484 ;
    END
  END w0_wd_in[195]
  PIN w0_wd_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 78.612 265.421 78.636 ;
    END
  END w0_wd_in[196]
  PIN w0_wd_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 79.764 265.421 79.788 ;
    END
  END w0_wd_in[197]
  PIN w0_wd_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 80.916 265.421 80.940 ;
    END
  END w0_wd_in[198]
  PIN w0_wd_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 82.068 265.421 82.092 ;
    END
  END w0_wd_in[199]
  PIN w0_wd_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 83.220 265.421 83.244 ;
    END
  END w0_wd_in[200]
  PIN w0_wd_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 84.372 265.421 84.396 ;
    END
  END w0_wd_in[201]
  PIN w0_wd_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 85.524 265.421 85.548 ;
    END
  END w0_wd_in[202]
  PIN w0_wd_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 86.676 265.421 86.700 ;
    END
  END w0_wd_in[203]
  PIN w0_wd_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 87.828 265.421 87.852 ;
    END
  END w0_wd_in[204]
  PIN w0_wd_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 88.980 265.421 89.004 ;
    END
  END w0_wd_in[205]
  PIN w0_wd_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 90.132 265.421 90.156 ;
    END
  END w0_wd_in[206]
  PIN w0_wd_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 91.284 265.421 91.308 ;
    END
  END w0_wd_in[207]
  PIN w0_wd_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 92.436 265.421 92.460 ;
    END
  END w0_wd_in[208]
  PIN w0_wd_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 93.588 265.421 93.612 ;
    END
  END w0_wd_in[209]
  PIN w0_wd_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 94.740 265.421 94.764 ;
    END
  END w0_wd_in[210]
  PIN w0_wd_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 95.892 265.421 95.916 ;
    END
  END w0_wd_in[211]
  PIN w0_wd_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 97.044 265.421 97.068 ;
    END
  END w0_wd_in[212]
  PIN w0_wd_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 98.196 265.421 98.220 ;
    END
  END w0_wd_in[213]
  PIN w0_wd_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 99.348 265.421 99.372 ;
    END
  END w0_wd_in[214]
  PIN w0_wd_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 100.500 265.421 100.524 ;
    END
  END w0_wd_in[215]
  PIN w0_wd_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 101.652 265.421 101.676 ;
    END
  END w0_wd_in[216]
  PIN w0_wd_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 102.804 265.421 102.828 ;
    END
  END w0_wd_in[217]
  PIN w0_wd_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 103.956 265.421 103.980 ;
    END
  END w0_wd_in[218]
  PIN w0_wd_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 105.108 265.421 105.132 ;
    END
  END w0_wd_in[219]
  PIN w0_wd_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 106.260 265.421 106.284 ;
    END
  END w0_wd_in[220]
  PIN w0_wd_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 107.412 265.421 107.436 ;
    END
  END w0_wd_in[221]
  PIN w0_wd_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 108.564 265.421 108.588 ;
    END
  END w0_wd_in[222]
  PIN w0_wd_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 109.716 265.421 109.740 ;
    END
  END w0_wd_in[223]
  PIN w0_wd_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 110.868 265.421 110.892 ;
    END
  END w0_wd_in[224]
  PIN w0_wd_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 112.020 265.421 112.044 ;
    END
  END w0_wd_in[225]
  PIN w0_wd_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 113.172 265.421 113.196 ;
    END
  END w0_wd_in[226]
  PIN w0_wd_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 114.324 265.421 114.348 ;
    END
  END w0_wd_in[227]
  PIN w0_wd_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 115.476 265.421 115.500 ;
    END
  END w0_wd_in[228]
  PIN w0_wd_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 116.628 265.421 116.652 ;
    END
  END w0_wd_in[229]
  PIN w0_wd_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 117.780 265.421 117.804 ;
    END
  END w0_wd_in[230]
  PIN w0_wd_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 118.932 265.421 118.956 ;
    END
  END w0_wd_in[231]
  PIN w0_wd_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 120.084 265.421 120.108 ;
    END
  END w0_wd_in[232]
  PIN w0_wd_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 121.236 265.421 121.260 ;
    END
  END w0_wd_in[233]
  PIN w0_wd_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 122.388 265.421 122.412 ;
    END
  END w0_wd_in[234]
  PIN w0_wd_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 123.540 265.421 123.564 ;
    END
  END w0_wd_in[235]
  PIN w0_wd_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 124.692 265.421 124.716 ;
    END
  END w0_wd_in[236]
  PIN w0_wd_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 125.844 265.421 125.868 ;
    END
  END w0_wd_in[237]
  PIN w0_wd_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 126.996 265.421 127.020 ;
    END
  END w0_wd_in[238]
  PIN w0_wd_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 128.148 265.421 128.172 ;
    END
  END w0_wd_in[239]
  PIN w0_wd_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 129.300 265.421 129.324 ;
    END
  END w0_wd_in[240]
  PIN w0_wd_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 130.452 265.421 130.476 ;
    END
  END w0_wd_in[241]
  PIN w0_wd_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 131.604 265.421 131.628 ;
    END
  END w0_wd_in[242]
  PIN w0_wd_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 132.756 265.421 132.780 ;
    END
  END w0_wd_in[243]
  PIN w0_wd_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 133.908 265.421 133.932 ;
    END
  END w0_wd_in[244]
  PIN w0_wd_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 135.060 265.421 135.084 ;
    END
  END w0_wd_in[245]
  PIN w0_wd_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 136.212 265.421 136.236 ;
    END
  END w0_wd_in[246]
  PIN w0_wd_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 137.364 265.421 137.388 ;
    END
  END w0_wd_in[247]
  PIN w0_wd_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 138.516 265.421 138.540 ;
    END
  END w0_wd_in[248]
  PIN w0_wd_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 139.668 265.421 139.692 ;
    END
  END w0_wd_in[249]
  PIN w0_wd_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 140.820 265.421 140.844 ;
    END
  END w0_wd_in[250]
  PIN w0_wd_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 141.972 265.421 141.996 ;
    END
  END w0_wd_in[251]
  PIN w0_wd_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 143.124 265.421 143.148 ;
    END
  END w0_wd_in[252]
  PIN w0_wd_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 144.276 265.421 144.300 ;
    END
  END w0_wd_in[253]
  PIN w0_wd_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 145.428 265.421 145.452 ;
    END
  END w0_wd_in[254]
  PIN w0_wd_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 146.580 265.421 146.604 ;
    END
  END w0_wd_in[255]
  PIN w0_wd_in[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 0.000 0.225 0.018 ;
    END
  END w0_wd_in[256]
  PIN w0_wd_in[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.711 0.000 0.729 0.018 ;
    END
  END w0_wd_in[257]
  PIN w0_wd_in[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.215 0.000 1.233 0.018 ;
    END
  END w0_wd_in[258]
  PIN w0_wd_in[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.719 0.000 1.737 0.018 ;
    END
  END w0_wd_in[259]
  PIN w0_wd_in[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.223 0.000 2.241 0.018 ;
    END
  END w0_wd_in[260]
  PIN w0_wd_in[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.727 0.000 2.745 0.018 ;
    END
  END w0_wd_in[261]
  PIN w0_wd_in[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.231 0.000 3.249 0.018 ;
    END
  END w0_wd_in[262]
  PIN w0_wd_in[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.735 0.000 3.753 0.018 ;
    END
  END w0_wd_in[263]
  PIN w0_wd_in[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.239 0.000 4.257 0.018 ;
    END
  END w0_wd_in[264]
  PIN w0_wd_in[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.743 0.000 4.761 0.018 ;
    END
  END w0_wd_in[265]
  PIN w0_wd_in[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.247 0.000 5.265 0.018 ;
    END
  END w0_wd_in[266]
  PIN w0_wd_in[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.751 0.000 5.769 0.018 ;
    END
  END w0_wd_in[267]
  PIN w0_wd_in[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.255 0.000 6.273 0.018 ;
    END
  END w0_wd_in[268]
  PIN w0_wd_in[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.759 0.000 6.777 0.018 ;
    END
  END w0_wd_in[269]
  PIN w0_wd_in[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.263 0.000 7.281 0.018 ;
    END
  END w0_wd_in[270]
  PIN w0_wd_in[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.767 0.000 7.785 0.018 ;
    END
  END w0_wd_in[271]
  PIN w0_wd_in[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.271 0.000 8.289 0.018 ;
    END
  END w0_wd_in[272]
  PIN w0_wd_in[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.775 0.000 8.793 0.018 ;
    END
  END w0_wd_in[273]
  PIN w0_wd_in[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.279 0.000 9.297 0.018 ;
    END
  END w0_wd_in[274]
  PIN w0_wd_in[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.783 0.000 9.801 0.018 ;
    END
  END w0_wd_in[275]
  PIN w0_wd_in[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.287 0.000 10.305 0.018 ;
    END
  END w0_wd_in[276]
  PIN w0_wd_in[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.791 0.000 10.809 0.018 ;
    END
  END w0_wd_in[277]
  PIN w0_wd_in[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 11.295 0.000 11.313 0.018 ;
    END
  END w0_wd_in[278]
  PIN w0_wd_in[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 11.799 0.000 11.817 0.018 ;
    END
  END w0_wd_in[279]
  PIN w0_wd_in[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.303 0.000 12.321 0.018 ;
    END
  END w0_wd_in[280]
  PIN w0_wd_in[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.807 0.000 12.825 0.018 ;
    END
  END w0_wd_in[281]
  PIN w0_wd_in[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 13.311 0.000 13.329 0.018 ;
    END
  END w0_wd_in[282]
  PIN w0_wd_in[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 13.815 0.000 13.833 0.018 ;
    END
  END w0_wd_in[283]
  PIN w0_wd_in[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 14.319 0.000 14.337 0.018 ;
    END
  END w0_wd_in[284]
  PIN w0_wd_in[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 14.823 0.000 14.841 0.018 ;
    END
  END w0_wd_in[285]
  PIN w0_wd_in[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 15.327 0.000 15.345 0.018 ;
    END
  END w0_wd_in[286]
  PIN w0_wd_in[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 15.831 0.000 15.849 0.018 ;
    END
  END w0_wd_in[287]
  PIN w0_wd_in[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 16.335 0.000 16.353 0.018 ;
    END
  END w0_wd_in[288]
  PIN w0_wd_in[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 16.839 0.000 16.857 0.018 ;
    END
  END w0_wd_in[289]
  PIN w0_wd_in[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 17.343 0.000 17.361 0.018 ;
    END
  END w0_wd_in[290]
  PIN w0_wd_in[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 17.847 0.000 17.865 0.018 ;
    END
  END w0_wd_in[291]
  PIN w0_wd_in[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 18.351 0.000 18.369 0.018 ;
    END
  END w0_wd_in[292]
  PIN w0_wd_in[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 18.855 0.000 18.873 0.018 ;
    END
  END w0_wd_in[293]
  PIN w0_wd_in[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 19.359 0.000 19.377 0.018 ;
    END
  END w0_wd_in[294]
  PIN w0_wd_in[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 19.863 0.000 19.881 0.018 ;
    END
  END w0_wd_in[295]
  PIN w0_wd_in[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 20.367 0.000 20.385 0.018 ;
    END
  END w0_wd_in[296]
  PIN w0_wd_in[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 20.871 0.000 20.889 0.018 ;
    END
  END w0_wd_in[297]
  PIN w0_wd_in[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 21.375 0.000 21.393 0.018 ;
    END
  END w0_wd_in[298]
  PIN w0_wd_in[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 21.879 0.000 21.897 0.018 ;
    END
  END w0_wd_in[299]
  PIN w0_wd_in[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 22.383 0.000 22.401 0.018 ;
    END
  END w0_wd_in[300]
  PIN w0_wd_in[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 22.887 0.000 22.905 0.018 ;
    END
  END w0_wd_in[301]
  PIN w0_wd_in[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 23.391 0.000 23.409 0.018 ;
    END
  END w0_wd_in[302]
  PIN w0_wd_in[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 23.895 0.000 23.913 0.018 ;
    END
  END w0_wd_in[303]
  PIN w0_wd_in[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 24.399 0.000 24.417 0.018 ;
    END
  END w0_wd_in[304]
  PIN w0_wd_in[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 24.903 0.000 24.921 0.018 ;
    END
  END w0_wd_in[305]
  PIN w0_wd_in[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 25.407 0.000 25.425 0.018 ;
    END
  END w0_wd_in[306]
  PIN w0_wd_in[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 25.911 0.000 25.929 0.018 ;
    END
  END w0_wd_in[307]
  PIN w0_wd_in[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 26.415 0.000 26.433 0.018 ;
    END
  END w0_wd_in[308]
  PIN w0_wd_in[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 26.919 0.000 26.937 0.018 ;
    END
  END w0_wd_in[309]
  PIN w0_wd_in[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 27.423 0.000 27.441 0.018 ;
    END
  END w0_wd_in[310]
  PIN w0_wd_in[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 27.927 0.000 27.945 0.018 ;
    END
  END w0_wd_in[311]
  PIN w0_wd_in[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 28.431 0.000 28.449 0.018 ;
    END
  END w0_wd_in[312]
  PIN w0_wd_in[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 28.935 0.000 28.953 0.018 ;
    END
  END w0_wd_in[313]
  PIN w0_wd_in[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 29.439 0.000 29.457 0.018 ;
    END
  END w0_wd_in[314]
  PIN w0_wd_in[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 29.943 0.000 29.961 0.018 ;
    END
  END w0_wd_in[315]
  PIN w0_wd_in[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 30.447 0.000 30.465 0.018 ;
    END
  END w0_wd_in[316]
  PIN w0_wd_in[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 30.951 0.000 30.969 0.018 ;
    END
  END w0_wd_in[317]
  PIN w0_wd_in[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 31.455 0.000 31.473 0.018 ;
    END
  END w0_wd_in[318]
  PIN w0_wd_in[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 31.959 0.000 31.977 0.018 ;
    END
  END w0_wd_in[319]
  PIN w0_wd_in[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 32.463 0.000 32.481 0.018 ;
    END
  END w0_wd_in[320]
  PIN w0_wd_in[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 32.967 0.000 32.985 0.018 ;
    END
  END w0_wd_in[321]
  PIN w0_wd_in[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 33.471 0.000 33.489 0.018 ;
    END
  END w0_wd_in[322]
  PIN w0_wd_in[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 33.975 0.000 33.993 0.018 ;
    END
  END w0_wd_in[323]
  PIN w0_wd_in[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 34.479 0.000 34.497 0.018 ;
    END
  END w0_wd_in[324]
  PIN w0_wd_in[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 34.983 0.000 35.001 0.018 ;
    END
  END w0_wd_in[325]
  PIN w0_wd_in[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 35.487 0.000 35.505 0.018 ;
    END
  END w0_wd_in[326]
  PIN w0_wd_in[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 35.991 0.000 36.009 0.018 ;
    END
  END w0_wd_in[327]
  PIN w0_wd_in[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 36.495 0.000 36.513 0.018 ;
    END
  END w0_wd_in[328]
  PIN w0_wd_in[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 36.999 0.000 37.017 0.018 ;
    END
  END w0_wd_in[329]
  PIN w0_wd_in[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 37.503 0.000 37.521 0.018 ;
    END
  END w0_wd_in[330]
  PIN w0_wd_in[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 38.007 0.000 38.025 0.018 ;
    END
  END w0_wd_in[331]
  PIN w0_wd_in[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 38.511 0.000 38.529 0.018 ;
    END
  END w0_wd_in[332]
  PIN w0_wd_in[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 39.015 0.000 39.033 0.018 ;
    END
  END w0_wd_in[333]
  PIN w0_wd_in[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 39.519 0.000 39.537 0.018 ;
    END
  END w0_wd_in[334]
  PIN w0_wd_in[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 40.023 0.000 40.041 0.018 ;
    END
  END w0_wd_in[335]
  PIN w0_wd_in[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 40.527 0.000 40.545 0.018 ;
    END
  END w0_wd_in[336]
  PIN w0_wd_in[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 41.031 0.000 41.049 0.018 ;
    END
  END w0_wd_in[337]
  PIN w0_wd_in[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 41.535 0.000 41.553 0.018 ;
    END
  END w0_wd_in[338]
  PIN w0_wd_in[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 42.039 0.000 42.057 0.018 ;
    END
  END w0_wd_in[339]
  PIN w0_wd_in[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 42.543 0.000 42.561 0.018 ;
    END
  END w0_wd_in[340]
  PIN w0_wd_in[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 43.047 0.000 43.065 0.018 ;
    END
  END w0_wd_in[341]
  PIN w0_wd_in[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 43.551 0.000 43.569 0.018 ;
    END
  END w0_wd_in[342]
  PIN w0_wd_in[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 44.055 0.000 44.073 0.018 ;
    END
  END w0_wd_in[343]
  PIN w0_wd_in[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 44.559 0.000 44.577 0.018 ;
    END
  END w0_wd_in[344]
  PIN w0_wd_in[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 45.063 0.000 45.081 0.018 ;
    END
  END w0_wd_in[345]
  PIN w0_wd_in[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 45.567 0.000 45.585 0.018 ;
    END
  END w0_wd_in[346]
  PIN w0_wd_in[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 46.071 0.000 46.089 0.018 ;
    END
  END w0_wd_in[347]
  PIN w0_wd_in[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 46.575 0.000 46.593 0.018 ;
    END
  END w0_wd_in[348]
  PIN w0_wd_in[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 47.079 0.000 47.097 0.018 ;
    END
  END w0_wd_in[349]
  PIN w0_wd_in[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 47.583 0.000 47.601 0.018 ;
    END
  END w0_wd_in[350]
  PIN w0_wd_in[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 48.087 0.000 48.105 0.018 ;
    END
  END w0_wd_in[351]
  PIN w0_wd_in[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 48.591 0.000 48.609 0.018 ;
    END
  END w0_wd_in[352]
  PIN w0_wd_in[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 49.095 0.000 49.113 0.018 ;
    END
  END w0_wd_in[353]
  PIN w0_wd_in[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 49.599 0.000 49.617 0.018 ;
    END
  END w0_wd_in[354]
  PIN w0_wd_in[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 50.103 0.000 50.121 0.018 ;
    END
  END w0_wd_in[355]
  PIN w0_wd_in[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 50.607 0.000 50.625 0.018 ;
    END
  END w0_wd_in[356]
  PIN w0_wd_in[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 51.111 0.000 51.129 0.018 ;
    END
  END w0_wd_in[357]
  PIN w0_wd_in[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 51.615 0.000 51.633 0.018 ;
    END
  END w0_wd_in[358]
  PIN w0_wd_in[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 52.119 0.000 52.137 0.018 ;
    END
  END w0_wd_in[359]
  PIN w0_wd_in[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 52.623 0.000 52.641 0.018 ;
    END
  END w0_wd_in[360]
  PIN w0_wd_in[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 53.127 0.000 53.145 0.018 ;
    END
  END w0_wd_in[361]
  PIN w0_wd_in[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 53.631 0.000 53.649 0.018 ;
    END
  END w0_wd_in[362]
  PIN w0_wd_in[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 54.135 0.000 54.153 0.018 ;
    END
  END w0_wd_in[363]
  PIN w0_wd_in[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 54.639 0.000 54.657 0.018 ;
    END
  END w0_wd_in[364]
  PIN w0_wd_in[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 55.143 0.000 55.161 0.018 ;
    END
  END w0_wd_in[365]
  PIN w0_wd_in[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 55.647 0.000 55.665 0.018 ;
    END
  END w0_wd_in[366]
  PIN w0_wd_in[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 56.151 0.000 56.169 0.018 ;
    END
  END w0_wd_in[367]
  PIN w0_wd_in[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 56.655 0.000 56.673 0.018 ;
    END
  END w0_wd_in[368]
  PIN w0_wd_in[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 57.159 0.000 57.177 0.018 ;
    END
  END w0_wd_in[369]
  PIN w0_wd_in[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 57.663 0.000 57.681 0.018 ;
    END
  END w0_wd_in[370]
  PIN w0_wd_in[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 58.167 0.000 58.185 0.018 ;
    END
  END w0_wd_in[371]
  PIN w0_wd_in[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 58.671 0.000 58.689 0.018 ;
    END
  END w0_wd_in[372]
  PIN w0_wd_in[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 59.175 0.000 59.193 0.018 ;
    END
  END w0_wd_in[373]
  PIN w0_wd_in[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 59.679 0.000 59.697 0.018 ;
    END
  END w0_wd_in[374]
  PIN w0_wd_in[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 60.183 0.000 60.201 0.018 ;
    END
  END w0_wd_in[375]
  PIN w0_wd_in[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 60.687 0.000 60.705 0.018 ;
    END
  END w0_wd_in[376]
  PIN w0_wd_in[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 61.191 0.000 61.209 0.018 ;
    END
  END w0_wd_in[377]
  PIN w0_wd_in[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 61.695 0.000 61.713 0.018 ;
    END
  END w0_wd_in[378]
  PIN w0_wd_in[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 62.199 0.000 62.217 0.018 ;
    END
  END w0_wd_in[379]
  PIN w0_wd_in[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 62.703 0.000 62.721 0.018 ;
    END
  END w0_wd_in[380]
  PIN w0_wd_in[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 63.207 0.000 63.225 0.018 ;
    END
  END w0_wd_in[381]
  PIN w0_wd_in[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 63.711 0.000 63.729 0.018 ;
    END
  END w0_wd_in[382]
  PIN w0_wd_in[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 64.215 0.000 64.233 0.018 ;
    END
  END w0_wd_in[383]
  PIN w0_wd_in[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 64.719 0.000 64.737 0.018 ;
    END
  END w0_wd_in[384]
  PIN w0_wd_in[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 65.223 0.000 65.241 0.018 ;
    END
  END w0_wd_in[385]
  PIN w0_wd_in[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 65.727 0.000 65.745 0.018 ;
    END
  END w0_wd_in[386]
  PIN w0_wd_in[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 66.231 0.000 66.249 0.018 ;
    END
  END w0_wd_in[387]
  PIN w0_wd_in[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 66.735 0.000 66.753 0.018 ;
    END
  END w0_wd_in[388]
  PIN w0_wd_in[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 67.239 0.000 67.257 0.018 ;
    END
  END w0_wd_in[389]
  PIN w0_wd_in[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 67.743 0.000 67.761 0.018 ;
    END
  END w0_wd_in[390]
  PIN w0_wd_in[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 68.247 0.000 68.265 0.018 ;
    END
  END w0_wd_in[391]
  PIN w0_wd_in[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 68.751 0.000 68.769 0.018 ;
    END
  END w0_wd_in[392]
  PIN w0_wd_in[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 69.255 0.000 69.273 0.018 ;
    END
  END w0_wd_in[393]
  PIN w0_wd_in[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 69.759 0.000 69.777 0.018 ;
    END
  END w0_wd_in[394]
  PIN w0_wd_in[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 70.263 0.000 70.281 0.018 ;
    END
  END w0_wd_in[395]
  PIN w0_wd_in[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 70.767 0.000 70.785 0.018 ;
    END
  END w0_wd_in[396]
  PIN w0_wd_in[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 71.271 0.000 71.289 0.018 ;
    END
  END w0_wd_in[397]
  PIN w0_wd_in[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 71.775 0.000 71.793 0.018 ;
    END
  END w0_wd_in[398]
  PIN w0_wd_in[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 72.279 0.000 72.297 0.018 ;
    END
  END w0_wd_in[399]
  PIN w0_wd_in[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 72.783 0.000 72.801 0.018 ;
    END
  END w0_wd_in[400]
  PIN w0_wd_in[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 73.287 0.000 73.305 0.018 ;
    END
  END w0_wd_in[401]
  PIN w0_wd_in[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 73.791 0.000 73.809 0.018 ;
    END
  END w0_wd_in[402]
  PIN w0_wd_in[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 74.295 0.000 74.313 0.018 ;
    END
  END w0_wd_in[403]
  PIN w0_wd_in[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 74.799 0.000 74.817 0.018 ;
    END
  END w0_wd_in[404]
  PIN w0_wd_in[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 75.303 0.000 75.321 0.018 ;
    END
  END w0_wd_in[405]
  PIN w0_wd_in[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 75.807 0.000 75.825 0.018 ;
    END
  END w0_wd_in[406]
  PIN w0_wd_in[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 76.311 0.000 76.329 0.018 ;
    END
  END w0_wd_in[407]
  PIN w0_wd_in[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 76.815 0.000 76.833 0.018 ;
    END
  END w0_wd_in[408]
  PIN w0_wd_in[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 77.319 0.000 77.337 0.018 ;
    END
  END w0_wd_in[409]
  PIN w0_wd_in[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 77.823 0.000 77.841 0.018 ;
    END
  END w0_wd_in[410]
  PIN w0_wd_in[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 78.327 0.000 78.345 0.018 ;
    END
  END w0_wd_in[411]
  PIN w0_wd_in[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 78.831 0.000 78.849 0.018 ;
    END
  END w0_wd_in[412]
  PIN w0_wd_in[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 79.335 0.000 79.353 0.018 ;
    END
  END w0_wd_in[413]
  PIN w0_wd_in[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 79.839 0.000 79.857 0.018 ;
    END
  END w0_wd_in[414]
  PIN w0_wd_in[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 80.343 0.000 80.361 0.018 ;
    END
  END w0_wd_in[415]
  PIN w0_wd_in[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 80.847 0.000 80.865 0.018 ;
    END
  END w0_wd_in[416]
  PIN w0_wd_in[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 81.351 0.000 81.369 0.018 ;
    END
  END w0_wd_in[417]
  PIN w0_wd_in[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 81.855 0.000 81.873 0.018 ;
    END
  END w0_wd_in[418]
  PIN w0_wd_in[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 82.359 0.000 82.377 0.018 ;
    END
  END w0_wd_in[419]
  PIN w0_wd_in[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 82.863 0.000 82.881 0.018 ;
    END
  END w0_wd_in[420]
  PIN w0_wd_in[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 83.367 0.000 83.385 0.018 ;
    END
  END w0_wd_in[421]
  PIN w0_wd_in[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 83.871 0.000 83.889 0.018 ;
    END
  END w0_wd_in[422]
  PIN w0_wd_in[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 84.375 0.000 84.393 0.018 ;
    END
  END w0_wd_in[423]
  PIN w0_wd_in[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 84.879 0.000 84.897 0.018 ;
    END
  END w0_wd_in[424]
  PIN w0_wd_in[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 85.383 0.000 85.401 0.018 ;
    END
  END w0_wd_in[425]
  PIN w0_wd_in[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 85.887 0.000 85.905 0.018 ;
    END
  END w0_wd_in[426]
  PIN w0_wd_in[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 86.391 0.000 86.409 0.018 ;
    END
  END w0_wd_in[427]
  PIN w0_wd_in[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 86.895 0.000 86.913 0.018 ;
    END
  END w0_wd_in[428]
  PIN w0_wd_in[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 87.399 0.000 87.417 0.018 ;
    END
  END w0_wd_in[429]
  PIN w0_wd_in[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 87.903 0.000 87.921 0.018 ;
    END
  END w0_wd_in[430]
  PIN w0_wd_in[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 88.407 0.000 88.425 0.018 ;
    END
  END w0_wd_in[431]
  PIN w0_wd_in[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 88.911 0.000 88.929 0.018 ;
    END
  END w0_wd_in[432]
  PIN w0_wd_in[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 89.415 0.000 89.433 0.018 ;
    END
  END w0_wd_in[433]
  PIN w0_wd_in[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 89.919 0.000 89.937 0.018 ;
    END
  END w0_wd_in[434]
  PIN w0_wd_in[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 90.423 0.000 90.441 0.018 ;
    END
  END w0_wd_in[435]
  PIN w0_wd_in[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 90.927 0.000 90.945 0.018 ;
    END
  END w0_wd_in[436]
  PIN w0_wd_in[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 91.431 0.000 91.449 0.018 ;
    END
  END w0_wd_in[437]
  PIN w0_wd_in[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 91.935 0.000 91.953 0.018 ;
    END
  END w0_wd_in[438]
  PIN w0_wd_in[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 92.439 0.000 92.457 0.018 ;
    END
  END w0_wd_in[439]
  PIN w0_wd_in[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 92.943 0.000 92.961 0.018 ;
    END
  END w0_wd_in[440]
  PIN w0_wd_in[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 93.447 0.000 93.465 0.018 ;
    END
  END w0_wd_in[441]
  PIN w0_wd_in[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 93.951 0.000 93.969 0.018 ;
    END
  END w0_wd_in[442]
  PIN w0_wd_in[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 94.455 0.000 94.473 0.018 ;
    END
  END w0_wd_in[443]
  PIN w0_wd_in[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 94.959 0.000 94.977 0.018 ;
    END
  END w0_wd_in[444]
  PIN w0_wd_in[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 95.463 0.000 95.481 0.018 ;
    END
  END w0_wd_in[445]
  PIN w0_wd_in[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 95.967 0.000 95.985 0.018 ;
    END
  END w0_wd_in[446]
  PIN w0_wd_in[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 96.471 0.000 96.489 0.018 ;
    END
  END w0_wd_in[447]
  PIN w0_wd_in[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 96.975 0.000 96.993 0.018 ;
    END
  END w0_wd_in[448]
  PIN w0_wd_in[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 97.479 0.000 97.497 0.018 ;
    END
  END w0_wd_in[449]
  PIN w0_wd_in[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 97.983 0.000 98.001 0.018 ;
    END
  END w0_wd_in[450]
  PIN w0_wd_in[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 98.487 0.000 98.505 0.018 ;
    END
  END w0_wd_in[451]
  PIN w0_wd_in[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 98.991 0.000 99.009 0.018 ;
    END
  END w0_wd_in[452]
  PIN w0_wd_in[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 99.495 0.000 99.513 0.018 ;
    END
  END w0_wd_in[453]
  PIN w0_wd_in[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 99.999 0.000 100.017 0.018 ;
    END
  END w0_wd_in[454]
  PIN w0_wd_in[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 100.503 0.000 100.521 0.018 ;
    END
  END w0_wd_in[455]
  PIN w0_wd_in[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 101.007 0.000 101.025 0.018 ;
    END
  END w0_wd_in[456]
  PIN w0_wd_in[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 101.511 0.000 101.529 0.018 ;
    END
  END w0_wd_in[457]
  PIN w0_wd_in[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 102.015 0.000 102.033 0.018 ;
    END
  END w0_wd_in[458]
  PIN w0_wd_in[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 102.519 0.000 102.537 0.018 ;
    END
  END w0_wd_in[459]
  PIN w0_wd_in[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 103.023 0.000 103.041 0.018 ;
    END
  END w0_wd_in[460]
  PIN w0_wd_in[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 103.527 0.000 103.545 0.018 ;
    END
  END w0_wd_in[461]
  PIN w0_wd_in[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 104.031 0.000 104.049 0.018 ;
    END
  END w0_wd_in[462]
  PIN w0_wd_in[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 104.535 0.000 104.553 0.018 ;
    END
  END w0_wd_in[463]
  PIN w0_wd_in[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 105.039 0.000 105.057 0.018 ;
    END
  END w0_wd_in[464]
  PIN w0_wd_in[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 105.543 0.000 105.561 0.018 ;
    END
  END w0_wd_in[465]
  PIN w0_wd_in[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 106.047 0.000 106.065 0.018 ;
    END
  END w0_wd_in[466]
  PIN w0_wd_in[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 106.551 0.000 106.569 0.018 ;
    END
  END w0_wd_in[467]
  PIN w0_wd_in[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 107.055 0.000 107.073 0.018 ;
    END
  END w0_wd_in[468]
  PIN w0_wd_in[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 107.559 0.000 107.577 0.018 ;
    END
  END w0_wd_in[469]
  PIN w0_wd_in[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 108.063 0.000 108.081 0.018 ;
    END
  END w0_wd_in[470]
  PIN w0_wd_in[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 108.567 0.000 108.585 0.018 ;
    END
  END w0_wd_in[471]
  PIN w0_wd_in[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 109.071 0.000 109.089 0.018 ;
    END
  END w0_wd_in[472]
  PIN w0_wd_in[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 109.575 0.000 109.593 0.018 ;
    END
  END w0_wd_in[473]
  PIN w0_wd_in[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 110.079 0.000 110.097 0.018 ;
    END
  END w0_wd_in[474]
  PIN w0_wd_in[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 110.583 0.000 110.601 0.018 ;
    END
  END w0_wd_in[475]
  PIN w0_wd_in[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 111.087 0.000 111.105 0.018 ;
    END
  END w0_wd_in[476]
  PIN w0_wd_in[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 111.591 0.000 111.609 0.018 ;
    END
  END w0_wd_in[477]
  PIN w0_wd_in[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 112.095 0.000 112.113 0.018 ;
    END
  END w0_wd_in[478]
  PIN w0_wd_in[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 112.599 0.000 112.617 0.018 ;
    END
  END w0_wd_in[479]
  PIN w0_wd_in[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 113.103 0.000 113.121 0.018 ;
    END
  END w0_wd_in[480]
  PIN w0_wd_in[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 113.607 0.000 113.625 0.018 ;
    END
  END w0_wd_in[481]
  PIN w0_wd_in[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 114.111 0.000 114.129 0.018 ;
    END
  END w0_wd_in[482]
  PIN w0_wd_in[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 114.615 0.000 114.633 0.018 ;
    END
  END w0_wd_in[483]
  PIN w0_wd_in[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 115.119 0.000 115.137 0.018 ;
    END
  END w0_wd_in[484]
  PIN w0_wd_in[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 115.623 0.000 115.641 0.018 ;
    END
  END w0_wd_in[485]
  PIN w0_wd_in[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 116.127 0.000 116.145 0.018 ;
    END
  END w0_wd_in[486]
  PIN w0_wd_in[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 116.631 0.000 116.649 0.018 ;
    END
  END w0_wd_in[487]
  PIN w0_wd_in[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 117.135 0.000 117.153 0.018 ;
    END
  END w0_wd_in[488]
  PIN w0_wd_in[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 117.639 0.000 117.657 0.018 ;
    END
  END w0_wd_in[489]
  PIN w0_wd_in[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 118.143 0.000 118.161 0.018 ;
    END
  END w0_wd_in[490]
  PIN w0_wd_in[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 118.647 0.000 118.665 0.018 ;
    END
  END w0_wd_in[491]
  PIN w0_wd_in[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 119.151 0.000 119.169 0.018 ;
    END
  END w0_wd_in[492]
  PIN w0_wd_in[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 119.655 0.000 119.673 0.018 ;
    END
  END w0_wd_in[493]
  PIN w0_wd_in[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 120.159 0.000 120.177 0.018 ;
    END
  END w0_wd_in[494]
  PIN w0_wd_in[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 120.663 0.000 120.681 0.018 ;
    END
  END w0_wd_in[495]
  PIN w0_wd_in[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 121.167 0.000 121.185 0.018 ;
    END
  END w0_wd_in[496]
  PIN w0_wd_in[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 121.671 0.000 121.689 0.018 ;
    END
  END w0_wd_in[497]
  PIN w0_wd_in[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 122.175 0.000 122.193 0.018 ;
    END
  END w0_wd_in[498]
  PIN w0_wd_in[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 122.679 0.000 122.697 0.018 ;
    END
  END w0_wd_in[499]
  PIN w0_wd_in[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 123.183 0.000 123.201 0.018 ;
    END
  END w0_wd_in[500]
  PIN w0_wd_in[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 123.687 0.000 123.705 0.018 ;
    END
  END w0_wd_in[501]
  PIN w0_wd_in[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 124.191 0.000 124.209 0.018 ;
    END
  END w0_wd_in[502]
  PIN w0_wd_in[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 124.695 0.000 124.713 0.018 ;
    END
  END w0_wd_in[503]
  PIN w0_wd_in[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 125.199 0.000 125.217 0.018 ;
    END
  END w0_wd_in[504]
  PIN w0_wd_in[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 125.703 0.000 125.721 0.018 ;
    END
  END w0_wd_in[505]
  PIN w0_wd_in[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 126.207 0.000 126.225 0.018 ;
    END
  END w0_wd_in[506]
  PIN w0_wd_in[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 126.711 0.000 126.729 0.018 ;
    END
  END w0_wd_in[507]
  PIN w0_wd_in[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 127.215 0.000 127.233 0.018 ;
    END
  END w0_wd_in[508]
  PIN w0_wd_in[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 127.719 0.000 127.737 0.018 ;
    END
  END w0_wd_in[509]
  PIN w0_wd_in[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 128.223 0.000 128.241 0.018 ;
    END
  END w0_wd_in[510]
  PIN w0_wd_in[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 128.727 0.000 128.745 0.018 ;
    END
  END w0_wd_in[511]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 129.231 0.000 129.249 0.018 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 129.735 0.000 129.753 0.018 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 130.239 0.000 130.257 0.018 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 130.743 0.000 130.761 0.018 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 131.247 0.000 131.265 0.018 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 131.751 0.000 131.769 0.018 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 132.255 0.000 132.273 0.018 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 132.759 0.000 132.777 0.018 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 133.263 0.000 133.281 0.018 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 133.767 0.000 133.785 0.018 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 134.271 0.000 134.289 0.018 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 134.775 0.000 134.793 0.018 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 135.279 0.000 135.297 0.018 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 135.783 0.000 135.801 0.018 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 136.287 0.000 136.305 0.018 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 136.791 0.000 136.809 0.018 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 137.295 0.000 137.313 0.018 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 137.799 0.000 137.817 0.018 ;
    END
  END r0_rd_out[17]
  PIN r0_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 138.303 0.000 138.321 0.018 ;
    END
  END r0_rd_out[18]
  PIN r0_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 138.807 0.000 138.825 0.018 ;
    END
  END r0_rd_out[19]
  PIN r0_rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 139.311 0.000 139.329 0.018 ;
    END
  END r0_rd_out[20]
  PIN r0_rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 139.815 0.000 139.833 0.018 ;
    END
  END r0_rd_out[21]
  PIN r0_rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 140.319 0.000 140.337 0.018 ;
    END
  END r0_rd_out[22]
  PIN r0_rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 140.823 0.000 140.841 0.018 ;
    END
  END r0_rd_out[23]
  PIN r0_rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 141.327 0.000 141.345 0.018 ;
    END
  END r0_rd_out[24]
  PIN r0_rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 141.831 0.000 141.849 0.018 ;
    END
  END r0_rd_out[25]
  PIN r0_rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 142.335 0.000 142.353 0.018 ;
    END
  END r0_rd_out[26]
  PIN r0_rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 142.839 0.000 142.857 0.018 ;
    END
  END r0_rd_out[27]
  PIN r0_rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 143.343 0.000 143.361 0.018 ;
    END
  END r0_rd_out[28]
  PIN r0_rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 143.847 0.000 143.865 0.018 ;
    END
  END r0_rd_out[29]
  PIN r0_rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 144.351 0.000 144.369 0.018 ;
    END
  END r0_rd_out[30]
  PIN r0_rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 144.855 0.000 144.873 0.018 ;
    END
  END r0_rd_out[31]
  PIN r0_rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 145.359 0.000 145.377 0.018 ;
    END
  END r0_rd_out[32]
  PIN r0_rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 145.863 0.000 145.881 0.018 ;
    END
  END r0_rd_out[33]
  PIN r0_rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 146.367 0.000 146.385 0.018 ;
    END
  END r0_rd_out[34]
  PIN r0_rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 146.871 0.000 146.889 0.018 ;
    END
  END r0_rd_out[35]
  PIN r0_rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 147.375 0.000 147.393 0.018 ;
    END
  END r0_rd_out[36]
  PIN r0_rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 147.879 0.000 147.897 0.018 ;
    END
  END r0_rd_out[37]
  PIN r0_rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 148.383 0.000 148.401 0.018 ;
    END
  END r0_rd_out[38]
  PIN r0_rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 148.887 0.000 148.905 0.018 ;
    END
  END r0_rd_out[39]
  PIN r0_rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 149.391 0.000 149.409 0.018 ;
    END
  END r0_rd_out[40]
  PIN r0_rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 149.895 0.000 149.913 0.018 ;
    END
  END r0_rd_out[41]
  PIN r0_rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 150.399 0.000 150.417 0.018 ;
    END
  END r0_rd_out[42]
  PIN r0_rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 150.903 0.000 150.921 0.018 ;
    END
  END r0_rd_out[43]
  PIN r0_rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 151.407 0.000 151.425 0.018 ;
    END
  END r0_rd_out[44]
  PIN r0_rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 151.911 0.000 151.929 0.018 ;
    END
  END r0_rd_out[45]
  PIN r0_rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 152.415 0.000 152.433 0.018 ;
    END
  END r0_rd_out[46]
  PIN r0_rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 152.919 0.000 152.937 0.018 ;
    END
  END r0_rd_out[47]
  PIN r0_rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 153.423 0.000 153.441 0.018 ;
    END
  END r0_rd_out[48]
  PIN r0_rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 153.927 0.000 153.945 0.018 ;
    END
  END r0_rd_out[49]
  PIN r0_rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 154.431 0.000 154.449 0.018 ;
    END
  END r0_rd_out[50]
  PIN r0_rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 154.935 0.000 154.953 0.018 ;
    END
  END r0_rd_out[51]
  PIN r0_rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 155.439 0.000 155.457 0.018 ;
    END
  END r0_rd_out[52]
  PIN r0_rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 155.943 0.000 155.961 0.018 ;
    END
  END r0_rd_out[53]
  PIN r0_rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 156.447 0.000 156.465 0.018 ;
    END
  END r0_rd_out[54]
  PIN r0_rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 156.951 0.000 156.969 0.018 ;
    END
  END r0_rd_out[55]
  PIN r0_rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 157.455 0.000 157.473 0.018 ;
    END
  END r0_rd_out[56]
  PIN r0_rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 157.959 0.000 157.977 0.018 ;
    END
  END r0_rd_out[57]
  PIN r0_rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 158.463 0.000 158.481 0.018 ;
    END
  END r0_rd_out[58]
  PIN r0_rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 158.967 0.000 158.985 0.018 ;
    END
  END r0_rd_out[59]
  PIN r0_rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 159.471 0.000 159.489 0.018 ;
    END
  END r0_rd_out[60]
  PIN r0_rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 159.975 0.000 159.993 0.018 ;
    END
  END r0_rd_out[61]
  PIN r0_rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 160.479 0.000 160.497 0.018 ;
    END
  END r0_rd_out[62]
  PIN r0_rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 160.983 0.000 161.001 0.018 ;
    END
  END r0_rd_out[63]
  PIN r0_rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 161.487 0.000 161.505 0.018 ;
    END
  END r0_rd_out[64]
  PIN r0_rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 161.991 0.000 162.009 0.018 ;
    END
  END r0_rd_out[65]
  PIN r0_rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 162.495 0.000 162.513 0.018 ;
    END
  END r0_rd_out[66]
  PIN r0_rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 162.999 0.000 163.017 0.018 ;
    END
  END r0_rd_out[67]
  PIN r0_rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 163.503 0.000 163.521 0.018 ;
    END
  END r0_rd_out[68]
  PIN r0_rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 164.007 0.000 164.025 0.018 ;
    END
  END r0_rd_out[69]
  PIN r0_rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 164.511 0.000 164.529 0.018 ;
    END
  END r0_rd_out[70]
  PIN r0_rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 165.015 0.000 165.033 0.018 ;
    END
  END r0_rd_out[71]
  PIN r0_rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 165.519 0.000 165.537 0.018 ;
    END
  END r0_rd_out[72]
  PIN r0_rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 166.023 0.000 166.041 0.018 ;
    END
  END r0_rd_out[73]
  PIN r0_rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 166.527 0.000 166.545 0.018 ;
    END
  END r0_rd_out[74]
  PIN r0_rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 167.031 0.000 167.049 0.018 ;
    END
  END r0_rd_out[75]
  PIN r0_rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 167.535 0.000 167.553 0.018 ;
    END
  END r0_rd_out[76]
  PIN r0_rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 168.039 0.000 168.057 0.018 ;
    END
  END r0_rd_out[77]
  PIN r0_rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 168.543 0.000 168.561 0.018 ;
    END
  END r0_rd_out[78]
  PIN r0_rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 169.047 0.000 169.065 0.018 ;
    END
  END r0_rd_out[79]
  PIN r0_rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 169.551 0.000 169.569 0.018 ;
    END
  END r0_rd_out[80]
  PIN r0_rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 170.055 0.000 170.073 0.018 ;
    END
  END r0_rd_out[81]
  PIN r0_rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 170.559 0.000 170.577 0.018 ;
    END
  END r0_rd_out[82]
  PIN r0_rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 171.063 0.000 171.081 0.018 ;
    END
  END r0_rd_out[83]
  PIN r0_rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 171.567 0.000 171.585 0.018 ;
    END
  END r0_rd_out[84]
  PIN r0_rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 172.071 0.000 172.089 0.018 ;
    END
  END r0_rd_out[85]
  PIN r0_rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 172.575 0.000 172.593 0.018 ;
    END
  END r0_rd_out[86]
  PIN r0_rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 173.079 0.000 173.097 0.018 ;
    END
  END r0_rd_out[87]
  PIN r0_rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 173.583 0.000 173.601 0.018 ;
    END
  END r0_rd_out[88]
  PIN r0_rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 174.087 0.000 174.105 0.018 ;
    END
  END r0_rd_out[89]
  PIN r0_rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 174.591 0.000 174.609 0.018 ;
    END
  END r0_rd_out[90]
  PIN r0_rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 175.095 0.000 175.113 0.018 ;
    END
  END r0_rd_out[91]
  PIN r0_rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 175.599 0.000 175.617 0.018 ;
    END
  END r0_rd_out[92]
  PIN r0_rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 176.103 0.000 176.121 0.018 ;
    END
  END r0_rd_out[93]
  PIN r0_rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 176.607 0.000 176.625 0.018 ;
    END
  END r0_rd_out[94]
  PIN r0_rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 177.111 0.000 177.129 0.018 ;
    END
  END r0_rd_out[95]
  PIN r0_rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 177.615 0.000 177.633 0.018 ;
    END
  END r0_rd_out[96]
  PIN r0_rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 178.119 0.000 178.137 0.018 ;
    END
  END r0_rd_out[97]
  PIN r0_rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 178.623 0.000 178.641 0.018 ;
    END
  END r0_rd_out[98]
  PIN r0_rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 179.127 0.000 179.145 0.018 ;
    END
  END r0_rd_out[99]
  PIN r0_rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 179.631 0.000 179.649 0.018 ;
    END
  END r0_rd_out[100]
  PIN r0_rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 180.135 0.000 180.153 0.018 ;
    END
  END r0_rd_out[101]
  PIN r0_rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 180.639 0.000 180.657 0.018 ;
    END
  END r0_rd_out[102]
  PIN r0_rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 181.143 0.000 181.161 0.018 ;
    END
  END r0_rd_out[103]
  PIN r0_rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 181.647 0.000 181.665 0.018 ;
    END
  END r0_rd_out[104]
  PIN r0_rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 182.151 0.000 182.169 0.018 ;
    END
  END r0_rd_out[105]
  PIN r0_rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 182.655 0.000 182.673 0.018 ;
    END
  END r0_rd_out[106]
  PIN r0_rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 183.159 0.000 183.177 0.018 ;
    END
  END r0_rd_out[107]
  PIN r0_rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 183.663 0.000 183.681 0.018 ;
    END
  END r0_rd_out[108]
  PIN r0_rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 184.167 0.000 184.185 0.018 ;
    END
  END r0_rd_out[109]
  PIN r0_rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 184.671 0.000 184.689 0.018 ;
    END
  END r0_rd_out[110]
  PIN r0_rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 185.175 0.000 185.193 0.018 ;
    END
  END r0_rd_out[111]
  PIN r0_rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 185.679 0.000 185.697 0.018 ;
    END
  END r0_rd_out[112]
  PIN r0_rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 186.183 0.000 186.201 0.018 ;
    END
  END r0_rd_out[113]
  PIN r0_rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 186.687 0.000 186.705 0.018 ;
    END
  END r0_rd_out[114]
  PIN r0_rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 187.191 0.000 187.209 0.018 ;
    END
  END r0_rd_out[115]
  PIN r0_rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 187.695 0.000 187.713 0.018 ;
    END
  END r0_rd_out[116]
  PIN r0_rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 188.199 0.000 188.217 0.018 ;
    END
  END r0_rd_out[117]
  PIN r0_rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 188.703 0.000 188.721 0.018 ;
    END
  END r0_rd_out[118]
  PIN r0_rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 189.207 0.000 189.225 0.018 ;
    END
  END r0_rd_out[119]
  PIN r0_rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 189.711 0.000 189.729 0.018 ;
    END
  END r0_rd_out[120]
  PIN r0_rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 190.215 0.000 190.233 0.018 ;
    END
  END r0_rd_out[121]
  PIN r0_rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 190.719 0.000 190.737 0.018 ;
    END
  END r0_rd_out[122]
  PIN r0_rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 191.223 0.000 191.241 0.018 ;
    END
  END r0_rd_out[123]
  PIN r0_rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 191.727 0.000 191.745 0.018 ;
    END
  END r0_rd_out[124]
  PIN r0_rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 192.231 0.000 192.249 0.018 ;
    END
  END r0_rd_out[125]
  PIN r0_rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 192.735 0.000 192.753 0.018 ;
    END
  END r0_rd_out[126]
  PIN r0_rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 193.239 0.000 193.257 0.018 ;
    END
  END r0_rd_out[127]
  PIN r0_rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 193.743 0.000 193.761 0.018 ;
    END
  END r0_rd_out[128]
  PIN r0_rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 194.247 0.000 194.265 0.018 ;
    END
  END r0_rd_out[129]
  PIN r0_rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 194.751 0.000 194.769 0.018 ;
    END
  END r0_rd_out[130]
  PIN r0_rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 195.255 0.000 195.273 0.018 ;
    END
  END r0_rd_out[131]
  PIN r0_rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 195.759 0.000 195.777 0.018 ;
    END
  END r0_rd_out[132]
  PIN r0_rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 196.263 0.000 196.281 0.018 ;
    END
  END r0_rd_out[133]
  PIN r0_rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 196.767 0.000 196.785 0.018 ;
    END
  END r0_rd_out[134]
  PIN r0_rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 197.271 0.000 197.289 0.018 ;
    END
  END r0_rd_out[135]
  PIN r0_rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 197.775 0.000 197.793 0.018 ;
    END
  END r0_rd_out[136]
  PIN r0_rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 198.279 0.000 198.297 0.018 ;
    END
  END r0_rd_out[137]
  PIN r0_rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 198.783 0.000 198.801 0.018 ;
    END
  END r0_rd_out[138]
  PIN r0_rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 199.287 0.000 199.305 0.018 ;
    END
  END r0_rd_out[139]
  PIN r0_rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 199.791 0.000 199.809 0.018 ;
    END
  END r0_rd_out[140]
  PIN r0_rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 200.295 0.000 200.313 0.018 ;
    END
  END r0_rd_out[141]
  PIN r0_rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 200.799 0.000 200.817 0.018 ;
    END
  END r0_rd_out[142]
  PIN r0_rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 201.303 0.000 201.321 0.018 ;
    END
  END r0_rd_out[143]
  PIN r0_rd_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 201.807 0.000 201.825 0.018 ;
    END
  END r0_rd_out[144]
  PIN r0_rd_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 202.311 0.000 202.329 0.018 ;
    END
  END r0_rd_out[145]
  PIN r0_rd_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 202.815 0.000 202.833 0.018 ;
    END
  END r0_rd_out[146]
  PIN r0_rd_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 203.319 0.000 203.337 0.018 ;
    END
  END r0_rd_out[147]
  PIN r0_rd_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 203.823 0.000 203.841 0.018 ;
    END
  END r0_rd_out[148]
  PIN r0_rd_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 204.327 0.000 204.345 0.018 ;
    END
  END r0_rd_out[149]
  PIN r0_rd_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 204.831 0.000 204.849 0.018 ;
    END
  END r0_rd_out[150]
  PIN r0_rd_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 205.335 0.000 205.353 0.018 ;
    END
  END r0_rd_out[151]
  PIN r0_rd_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 205.839 0.000 205.857 0.018 ;
    END
  END r0_rd_out[152]
  PIN r0_rd_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 206.343 0.000 206.361 0.018 ;
    END
  END r0_rd_out[153]
  PIN r0_rd_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 206.847 0.000 206.865 0.018 ;
    END
  END r0_rd_out[154]
  PIN r0_rd_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 207.351 0.000 207.369 0.018 ;
    END
  END r0_rd_out[155]
  PIN r0_rd_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 207.855 0.000 207.873 0.018 ;
    END
  END r0_rd_out[156]
  PIN r0_rd_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 208.359 0.000 208.377 0.018 ;
    END
  END r0_rd_out[157]
  PIN r0_rd_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 208.863 0.000 208.881 0.018 ;
    END
  END r0_rd_out[158]
  PIN r0_rd_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 209.367 0.000 209.385 0.018 ;
    END
  END r0_rd_out[159]
  PIN r0_rd_out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 209.871 0.000 209.889 0.018 ;
    END
  END r0_rd_out[160]
  PIN r0_rd_out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 210.375 0.000 210.393 0.018 ;
    END
  END r0_rd_out[161]
  PIN r0_rd_out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 210.879 0.000 210.897 0.018 ;
    END
  END r0_rd_out[162]
  PIN r0_rd_out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 211.383 0.000 211.401 0.018 ;
    END
  END r0_rd_out[163]
  PIN r0_rd_out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 211.887 0.000 211.905 0.018 ;
    END
  END r0_rd_out[164]
  PIN r0_rd_out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 212.391 0.000 212.409 0.018 ;
    END
  END r0_rd_out[165]
  PIN r0_rd_out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 212.895 0.000 212.913 0.018 ;
    END
  END r0_rd_out[166]
  PIN r0_rd_out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 213.399 0.000 213.417 0.018 ;
    END
  END r0_rd_out[167]
  PIN r0_rd_out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 213.903 0.000 213.921 0.018 ;
    END
  END r0_rd_out[168]
  PIN r0_rd_out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 214.407 0.000 214.425 0.018 ;
    END
  END r0_rd_out[169]
  PIN r0_rd_out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 214.911 0.000 214.929 0.018 ;
    END
  END r0_rd_out[170]
  PIN r0_rd_out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 215.415 0.000 215.433 0.018 ;
    END
  END r0_rd_out[171]
  PIN r0_rd_out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 215.919 0.000 215.937 0.018 ;
    END
  END r0_rd_out[172]
  PIN r0_rd_out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 216.423 0.000 216.441 0.018 ;
    END
  END r0_rd_out[173]
  PIN r0_rd_out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 216.927 0.000 216.945 0.018 ;
    END
  END r0_rd_out[174]
  PIN r0_rd_out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 217.431 0.000 217.449 0.018 ;
    END
  END r0_rd_out[175]
  PIN r0_rd_out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 217.935 0.000 217.953 0.018 ;
    END
  END r0_rd_out[176]
  PIN r0_rd_out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 218.439 0.000 218.457 0.018 ;
    END
  END r0_rd_out[177]
  PIN r0_rd_out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 218.943 0.000 218.961 0.018 ;
    END
  END r0_rd_out[178]
  PIN r0_rd_out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 219.447 0.000 219.465 0.018 ;
    END
  END r0_rd_out[179]
  PIN r0_rd_out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 219.951 0.000 219.969 0.018 ;
    END
  END r0_rd_out[180]
  PIN r0_rd_out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 220.455 0.000 220.473 0.018 ;
    END
  END r0_rd_out[181]
  PIN r0_rd_out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 220.959 0.000 220.977 0.018 ;
    END
  END r0_rd_out[182]
  PIN r0_rd_out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 221.463 0.000 221.481 0.018 ;
    END
  END r0_rd_out[183]
  PIN r0_rd_out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 221.967 0.000 221.985 0.018 ;
    END
  END r0_rd_out[184]
  PIN r0_rd_out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 222.471 0.000 222.489 0.018 ;
    END
  END r0_rd_out[185]
  PIN r0_rd_out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 222.975 0.000 222.993 0.018 ;
    END
  END r0_rd_out[186]
  PIN r0_rd_out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 223.479 0.000 223.497 0.018 ;
    END
  END r0_rd_out[187]
  PIN r0_rd_out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 223.983 0.000 224.001 0.018 ;
    END
  END r0_rd_out[188]
  PIN r0_rd_out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 224.487 0.000 224.505 0.018 ;
    END
  END r0_rd_out[189]
  PIN r0_rd_out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 224.991 0.000 225.009 0.018 ;
    END
  END r0_rd_out[190]
  PIN r0_rd_out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 225.495 0.000 225.513 0.018 ;
    END
  END r0_rd_out[191]
  PIN r0_rd_out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 225.999 0.000 226.017 0.018 ;
    END
  END r0_rd_out[192]
  PIN r0_rd_out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 226.503 0.000 226.521 0.018 ;
    END
  END r0_rd_out[193]
  PIN r0_rd_out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 227.007 0.000 227.025 0.018 ;
    END
  END r0_rd_out[194]
  PIN r0_rd_out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 227.511 0.000 227.529 0.018 ;
    END
  END r0_rd_out[195]
  PIN r0_rd_out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 228.015 0.000 228.033 0.018 ;
    END
  END r0_rd_out[196]
  PIN r0_rd_out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 228.519 0.000 228.537 0.018 ;
    END
  END r0_rd_out[197]
  PIN r0_rd_out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 229.023 0.000 229.041 0.018 ;
    END
  END r0_rd_out[198]
  PIN r0_rd_out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 229.527 0.000 229.545 0.018 ;
    END
  END r0_rd_out[199]
  PIN r0_rd_out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 230.031 0.000 230.049 0.018 ;
    END
  END r0_rd_out[200]
  PIN r0_rd_out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 230.535 0.000 230.553 0.018 ;
    END
  END r0_rd_out[201]
  PIN r0_rd_out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 231.039 0.000 231.057 0.018 ;
    END
  END r0_rd_out[202]
  PIN r0_rd_out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 231.543 0.000 231.561 0.018 ;
    END
  END r0_rd_out[203]
  PIN r0_rd_out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 232.047 0.000 232.065 0.018 ;
    END
  END r0_rd_out[204]
  PIN r0_rd_out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 232.551 0.000 232.569 0.018 ;
    END
  END r0_rd_out[205]
  PIN r0_rd_out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 233.055 0.000 233.073 0.018 ;
    END
  END r0_rd_out[206]
  PIN r0_rd_out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 233.559 0.000 233.577 0.018 ;
    END
  END r0_rd_out[207]
  PIN r0_rd_out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 234.063 0.000 234.081 0.018 ;
    END
  END r0_rd_out[208]
  PIN r0_rd_out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 234.567 0.000 234.585 0.018 ;
    END
  END r0_rd_out[209]
  PIN r0_rd_out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 235.071 0.000 235.089 0.018 ;
    END
  END r0_rd_out[210]
  PIN r0_rd_out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 235.575 0.000 235.593 0.018 ;
    END
  END r0_rd_out[211]
  PIN r0_rd_out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 236.079 0.000 236.097 0.018 ;
    END
  END r0_rd_out[212]
  PIN r0_rd_out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 236.583 0.000 236.601 0.018 ;
    END
  END r0_rd_out[213]
  PIN r0_rd_out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 237.087 0.000 237.105 0.018 ;
    END
  END r0_rd_out[214]
  PIN r0_rd_out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 237.591 0.000 237.609 0.018 ;
    END
  END r0_rd_out[215]
  PIN r0_rd_out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 238.095 0.000 238.113 0.018 ;
    END
  END r0_rd_out[216]
  PIN r0_rd_out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 238.599 0.000 238.617 0.018 ;
    END
  END r0_rd_out[217]
  PIN r0_rd_out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 239.103 0.000 239.121 0.018 ;
    END
  END r0_rd_out[218]
  PIN r0_rd_out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 239.607 0.000 239.625 0.018 ;
    END
  END r0_rd_out[219]
  PIN r0_rd_out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 240.111 0.000 240.129 0.018 ;
    END
  END r0_rd_out[220]
  PIN r0_rd_out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 240.615 0.000 240.633 0.018 ;
    END
  END r0_rd_out[221]
  PIN r0_rd_out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 241.119 0.000 241.137 0.018 ;
    END
  END r0_rd_out[222]
  PIN r0_rd_out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 241.623 0.000 241.641 0.018 ;
    END
  END r0_rd_out[223]
  PIN r0_rd_out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 242.127 0.000 242.145 0.018 ;
    END
  END r0_rd_out[224]
  PIN r0_rd_out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 242.631 0.000 242.649 0.018 ;
    END
  END r0_rd_out[225]
  PIN r0_rd_out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 243.135 0.000 243.153 0.018 ;
    END
  END r0_rd_out[226]
  PIN r0_rd_out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 243.639 0.000 243.657 0.018 ;
    END
  END r0_rd_out[227]
  PIN r0_rd_out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 244.143 0.000 244.161 0.018 ;
    END
  END r0_rd_out[228]
  PIN r0_rd_out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 244.647 0.000 244.665 0.018 ;
    END
  END r0_rd_out[229]
  PIN r0_rd_out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 245.151 0.000 245.169 0.018 ;
    END
  END r0_rd_out[230]
  PIN r0_rd_out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 245.655 0.000 245.673 0.018 ;
    END
  END r0_rd_out[231]
  PIN r0_rd_out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 246.159 0.000 246.177 0.018 ;
    END
  END r0_rd_out[232]
  PIN r0_rd_out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 246.663 0.000 246.681 0.018 ;
    END
  END r0_rd_out[233]
  PIN r0_rd_out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 247.167 0.000 247.185 0.018 ;
    END
  END r0_rd_out[234]
  PIN r0_rd_out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 247.671 0.000 247.689 0.018 ;
    END
  END r0_rd_out[235]
  PIN r0_rd_out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 248.175 0.000 248.193 0.018 ;
    END
  END r0_rd_out[236]
  PIN r0_rd_out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 248.679 0.000 248.697 0.018 ;
    END
  END r0_rd_out[237]
  PIN r0_rd_out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 249.183 0.000 249.201 0.018 ;
    END
  END r0_rd_out[238]
  PIN r0_rd_out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 249.687 0.000 249.705 0.018 ;
    END
  END r0_rd_out[239]
  PIN r0_rd_out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 250.191 0.000 250.209 0.018 ;
    END
  END r0_rd_out[240]
  PIN r0_rd_out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 250.695 0.000 250.713 0.018 ;
    END
  END r0_rd_out[241]
  PIN r0_rd_out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 251.199 0.000 251.217 0.018 ;
    END
  END r0_rd_out[242]
  PIN r0_rd_out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 251.703 0.000 251.721 0.018 ;
    END
  END r0_rd_out[243]
  PIN r0_rd_out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 252.207 0.000 252.225 0.018 ;
    END
  END r0_rd_out[244]
  PIN r0_rd_out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 252.711 0.000 252.729 0.018 ;
    END
  END r0_rd_out[245]
  PIN r0_rd_out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 253.215 0.000 253.233 0.018 ;
    END
  END r0_rd_out[246]
  PIN r0_rd_out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 253.719 0.000 253.737 0.018 ;
    END
  END r0_rd_out[247]
  PIN r0_rd_out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 254.223 0.000 254.241 0.018 ;
    END
  END r0_rd_out[248]
  PIN r0_rd_out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 254.727 0.000 254.745 0.018 ;
    END
  END r0_rd_out[249]
  PIN r0_rd_out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 255.231 0.000 255.249 0.018 ;
    END
  END r0_rd_out[250]
  PIN r0_rd_out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 255.735 0.000 255.753 0.018 ;
    END
  END r0_rd_out[251]
  PIN r0_rd_out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 256.239 0.000 256.257 0.018 ;
    END
  END r0_rd_out[252]
  PIN r0_rd_out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 256.743 0.000 256.761 0.018 ;
    END
  END r0_rd_out[253]
  PIN r0_rd_out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 257.247 0.000 257.265 0.018 ;
    END
  END r0_rd_out[254]
  PIN r0_rd_out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 257.751 0.000 257.769 0.018 ;
    END
  END r0_rd_out[255]
  PIN r0_rd_out[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 165.870 0.225 165.888 ;
    END
  END r0_rd_out[256]
  PIN r0_rd_out[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.215 165.870 1.233 165.888 ;
    END
  END r0_rd_out[257]
  PIN r0_rd_out[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.223 165.870 2.241 165.888 ;
    END
  END r0_rd_out[258]
  PIN r0_rd_out[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.231 165.870 3.249 165.888 ;
    END
  END r0_rd_out[259]
  PIN r0_rd_out[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.239 165.870 4.257 165.888 ;
    END
  END r0_rd_out[260]
  PIN r0_rd_out[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.247 165.870 5.265 165.888 ;
    END
  END r0_rd_out[261]
  PIN r0_rd_out[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.255 165.870 6.273 165.888 ;
    END
  END r0_rd_out[262]
  PIN r0_rd_out[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.263 165.870 7.281 165.888 ;
    END
  END r0_rd_out[263]
  PIN r0_rd_out[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.271 165.870 8.289 165.888 ;
    END
  END r0_rd_out[264]
  PIN r0_rd_out[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.279 165.870 9.297 165.888 ;
    END
  END r0_rd_out[265]
  PIN r0_rd_out[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.287 165.870 10.305 165.888 ;
    END
  END r0_rd_out[266]
  PIN r0_rd_out[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 11.295 165.870 11.313 165.888 ;
    END
  END r0_rd_out[267]
  PIN r0_rd_out[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.303 165.870 12.321 165.888 ;
    END
  END r0_rd_out[268]
  PIN r0_rd_out[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 13.311 165.870 13.329 165.888 ;
    END
  END r0_rd_out[269]
  PIN r0_rd_out[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 14.319 165.870 14.337 165.888 ;
    END
  END r0_rd_out[270]
  PIN r0_rd_out[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 15.327 165.870 15.345 165.888 ;
    END
  END r0_rd_out[271]
  PIN r0_rd_out[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 16.335 165.870 16.353 165.888 ;
    END
  END r0_rd_out[272]
  PIN r0_rd_out[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 17.343 165.870 17.361 165.888 ;
    END
  END r0_rd_out[273]
  PIN r0_rd_out[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 18.351 165.870 18.369 165.888 ;
    END
  END r0_rd_out[274]
  PIN r0_rd_out[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 19.359 165.870 19.377 165.888 ;
    END
  END r0_rd_out[275]
  PIN r0_rd_out[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 20.367 165.870 20.385 165.888 ;
    END
  END r0_rd_out[276]
  PIN r0_rd_out[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 21.375 165.870 21.393 165.888 ;
    END
  END r0_rd_out[277]
  PIN r0_rd_out[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 22.383 165.870 22.401 165.888 ;
    END
  END r0_rd_out[278]
  PIN r0_rd_out[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 23.391 165.870 23.409 165.888 ;
    END
  END r0_rd_out[279]
  PIN r0_rd_out[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 24.399 165.870 24.417 165.888 ;
    END
  END r0_rd_out[280]
  PIN r0_rd_out[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 25.407 165.870 25.425 165.888 ;
    END
  END r0_rd_out[281]
  PIN r0_rd_out[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 26.415 165.870 26.433 165.888 ;
    END
  END r0_rd_out[282]
  PIN r0_rd_out[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 27.423 165.870 27.441 165.888 ;
    END
  END r0_rd_out[283]
  PIN r0_rd_out[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 28.431 165.870 28.449 165.888 ;
    END
  END r0_rd_out[284]
  PIN r0_rd_out[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 29.439 165.870 29.457 165.888 ;
    END
  END r0_rd_out[285]
  PIN r0_rd_out[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 30.447 165.870 30.465 165.888 ;
    END
  END r0_rd_out[286]
  PIN r0_rd_out[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 31.455 165.870 31.473 165.888 ;
    END
  END r0_rd_out[287]
  PIN r0_rd_out[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 32.463 165.870 32.481 165.888 ;
    END
  END r0_rd_out[288]
  PIN r0_rd_out[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 33.471 165.870 33.489 165.888 ;
    END
  END r0_rd_out[289]
  PIN r0_rd_out[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 34.479 165.870 34.497 165.888 ;
    END
  END r0_rd_out[290]
  PIN r0_rd_out[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 35.487 165.870 35.505 165.888 ;
    END
  END r0_rd_out[291]
  PIN r0_rd_out[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 36.495 165.870 36.513 165.888 ;
    END
  END r0_rd_out[292]
  PIN r0_rd_out[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 37.503 165.870 37.521 165.888 ;
    END
  END r0_rd_out[293]
  PIN r0_rd_out[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 38.511 165.870 38.529 165.888 ;
    END
  END r0_rd_out[294]
  PIN r0_rd_out[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 39.519 165.870 39.537 165.888 ;
    END
  END r0_rd_out[295]
  PIN r0_rd_out[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 40.527 165.870 40.545 165.888 ;
    END
  END r0_rd_out[296]
  PIN r0_rd_out[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 41.535 165.870 41.553 165.888 ;
    END
  END r0_rd_out[297]
  PIN r0_rd_out[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 42.543 165.870 42.561 165.888 ;
    END
  END r0_rd_out[298]
  PIN r0_rd_out[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 43.551 165.870 43.569 165.888 ;
    END
  END r0_rd_out[299]
  PIN r0_rd_out[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 44.559 165.870 44.577 165.888 ;
    END
  END r0_rd_out[300]
  PIN r0_rd_out[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 45.567 165.870 45.585 165.888 ;
    END
  END r0_rd_out[301]
  PIN r0_rd_out[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 46.575 165.870 46.593 165.888 ;
    END
  END r0_rd_out[302]
  PIN r0_rd_out[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 47.583 165.870 47.601 165.888 ;
    END
  END r0_rd_out[303]
  PIN r0_rd_out[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 48.591 165.870 48.609 165.888 ;
    END
  END r0_rd_out[304]
  PIN r0_rd_out[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 49.599 165.870 49.617 165.888 ;
    END
  END r0_rd_out[305]
  PIN r0_rd_out[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 50.607 165.870 50.625 165.888 ;
    END
  END r0_rd_out[306]
  PIN r0_rd_out[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 51.615 165.870 51.633 165.888 ;
    END
  END r0_rd_out[307]
  PIN r0_rd_out[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 52.623 165.870 52.641 165.888 ;
    END
  END r0_rd_out[308]
  PIN r0_rd_out[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 53.631 165.870 53.649 165.888 ;
    END
  END r0_rd_out[309]
  PIN r0_rd_out[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 54.639 165.870 54.657 165.888 ;
    END
  END r0_rd_out[310]
  PIN r0_rd_out[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 55.647 165.870 55.665 165.888 ;
    END
  END r0_rd_out[311]
  PIN r0_rd_out[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 56.655 165.870 56.673 165.888 ;
    END
  END r0_rd_out[312]
  PIN r0_rd_out[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 57.663 165.870 57.681 165.888 ;
    END
  END r0_rd_out[313]
  PIN r0_rd_out[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 58.671 165.870 58.689 165.888 ;
    END
  END r0_rd_out[314]
  PIN r0_rd_out[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 59.679 165.870 59.697 165.888 ;
    END
  END r0_rd_out[315]
  PIN r0_rd_out[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 60.687 165.870 60.705 165.888 ;
    END
  END r0_rd_out[316]
  PIN r0_rd_out[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 61.695 165.870 61.713 165.888 ;
    END
  END r0_rd_out[317]
  PIN r0_rd_out[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 62.703 165.870 62.721 165.888 ;
    END
  END r0_rd_out[318]
  PIN r0_rd_out[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 63.711 165.870 63.729 165.888 ;
    END
  END r0_rd_out[319]
  PIN r0_rd_out[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 64.719 165.870 64.737 165.888 ;
    END
  END r0_rd_out[320]
  PIN r0_rd_out[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 65.727 165.870 65.745 165.888 ;
    END
  END r0_rd_out[321]
  PIN r0_rd_out[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 66.735 165.870 66.753 165.888 ;
    END
  END r0_rd_out[322]
  PIN r0_rd_out[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 67.743 165.870 67.761 165.888 ;
    END
  END r0_rd_out[323]
  PIN r0_rd_out[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 68.751 165.870 68.769 165.888 ;
    END
  END r0_rd_out[324]
  PIN r0_rd_out[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 69.759 165.870 69.777 165.888 ;
    END
  END r0_rd_out[325]
  PIN r0_rd_out[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 70.767 165.870 70.785 165.888 ;
    END
  END r0_rd_out[326]
  PIN r0_rd_out[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 71.775 165.870 71.793 165.888 ;
    END
  END r0_rd_out[327]
  PIN r0_rd_out[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 72.783 165.870 72.801 165.888 ;
    END
  END r0_rd_out[328]
  PIN r0_rd_out[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 73.791 165.870 73.809 165.888 ;
    END
  END r0_rd_out[329]
  PIN r0_rd_out[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 74.799 165.870 74.817 165.888 ;
    END
  END r0_rd_out[330]
  PIN r0_rd_out[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 75.807 165.870 75.825 165.888 ;
    END
  END r0_rd_out[331]
  PIN r0_rd_out[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 76.815 165.870 76.833 165.888 ;
    END
  END r0_rd_out[332]
  PIN r0_rd_out[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 77.823 165.870 77.841 165.888 ;
    END
  END r0_rd_out[333]
  PIN r0_rd_out[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 78.831 165.870 78.849 165.888 ;
    END
  END r0_rd_out[334]
  PIN r0_rd_out[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 79.839 165.870 79.857 165.888 ;
    END
  END r0_rd_out[335]
  PIN r0_rd_out[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 80.847 165.870 80.865 165.888 ;
    END
  END r0_rd_out[336]
  PIN r0_rd_out[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 81.855 165.870 81.873 165.888 ;
    END
  END r0_rd_out[337]
  PIN r0_rd_out[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 82.863 165.870 82.881 165.888 ;
    END
  END r0_rd_out[338]
  PIN r0_rd_out[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 83.871 165.870 83.889 165.888 ;
    END
  END r0_rd_out[339]
  PIN r0_rd_out[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 84.879 165.870 84.897 165.888 ;
    END
  END r0_rd_out[340]
  PIN r0_rd_out[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 85.887 165.870 85.905 165.888 ;
    END
  END r0_rd_out[341]
  PIN r0_rd_out[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 86.895 165.870 86.913 165.888 ;
    END
  END r0_rd_out[342]
  PIN r0_rd_out[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 87.903 165.870 87.921 165.888 ;
    END
  END r0_rd_out[343]
  PIN r0_rd_out[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 88.911 165.870 88.929 165.888 ;
    END
  END r0_rd_out[344]
  PIN r0_rd_out[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 89.919 165.870 89.937 165.888 ;
    END
  END r0_rd_out[345]
  PIN r0_rd_out[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 90.927 165.870 90.945 165.888 ;
    END
  END r0_rd_out[346]
  PIN r0_rd_out[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 91.935 165.870 91.953 165.888 ;
    END
  END r0_rd_out[347]
  PIN r0_rd_out[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 92.943 165.870 92.961 165.888 ;
    END
  END r0_rd_out[348]
  PIN r0_rd_out[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 93.951 165.870 93.969 165.888 ;
    END
  END r0_rd_out[349]
  PIN r0_rd_out[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 94.959 165.870 94.977 165.888 ;
    END
  END r0_rd_out[350]
  PIN r0_rd_out[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 95.967 165.870 95.985 165.888 ;
    END
  END r0_rd_out[351]
  PIN r0_rd_out[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 96.975 165.870 96.993 165.888 ;
    END
  END r0_rd_out[352]
  PIN r0_rd_out[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 97.983 165.870 98.001 165.888 ;
    END
  END r0_rd_out[353]
  PIN r0_rd_out[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 98.991 165.870 99.009 165.888 ;
    END
  END r0_rd_out[354]
  PIN r0_rd_out[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 99.999 165.870 100.017 165.888 ;
    END
  END r0_rd_out[355]
  PIN r0_rd_out[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 101.007 165.870 101.025 165.888 ;
    END
  END r0_rd_out[356]
  PIN r0_rd_out[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 102.015 165.870 102.033 165.888 ;
    END
  END r0_rd_out[357]
  PIN r0_rd_out[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 103.023 165.870 103.041 165.888 ;
    END
  END r0_rd_out[358]
  PIN r0_rd_out[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 104.031 165.870 104.049 165.888 ;
    END
  END r0_rd_out[359]
  PIN r0_rd_out[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 105.039 165.870 105.057 165.888 ;
    END
  END r0_rd_out[360]
  PIN r0_rd_out[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 106.047 165.870 106.065 165.888 ;
    END
  END r0_rd_out[361]
  PIN r0_rd_out[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 107.055 165.870 107.073 165.888 ;
    END
  END r0_rd_out[362]
  PIN r0_rd_out[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 108.063 165.870 108.081 165.888 ;
    END
  END r0_rd_out[363]
  PIN r0_rd_out[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 109.071 165.870 109.089 165.888 ;
    END
  END r0_rd_out[364]
  PIN r0_rd_out[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 110.079 165.870 110.097 165.888 ;
    END
  END r0_rd_out[365]
  PIN r0_rd_out[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 111.087 165.870 111.105 165.888 ;
    END
  END r0_rd_out[366]
  PIN r0_rd_out[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 112.095 165.870 112.113 165.888 ;
    END
  END r0_rd_out[367]
  PIN r0_rd_out[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 113.103 165.870 113.121 165.888 ;
    END
  END r0_rd_out[368]
  PIN r0_rd_out[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 114.111 165.870 114.129 165.888 ;
    END
  END r0_rd_out[369]
  PIN r0_rd_out[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 115.119 165.870 115.137 165.888 ;
    END
  END r0_rd_out[370]
  PIN r0_rd_out[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 116.127 165.870 116.145 165.888 ;
    END
  END r0_rd_out[371]
  PIN r0_rd_out[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 117.135 165.870 117.153 165.888 ;
    END
  END r0_rd_out[372]
  PIN r0_rd_out[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 118.143 165.870 118.161 165.888 ;
    END
  END r0_rd_out[373]
  PIN r0_rd_out[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 119.151 165.870 119.169 165.888 ;
    END
  END r0_rd_out[374]
  PIN r0_rd_out[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 120.159 165.870 120.177 165.888 ;
    END
  END r0_rd_out[375]
  PIN r0_rd_out[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 121.167 165.870 121.185 165.888 ;
    END
  END r0_rd_out[376]
  PIN r0_rd_out[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 122.175 165.870 122.193 165.888 ;
    END
  END r0_rd_out[377]
  PIN r0_rd_out[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 123.183 165.870 123.201 165.888 ;
    END
  END r0_rd_out[378]
  PIN r0_rd_out[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 124.191 165.870 124.209 165.888 ;
    END
  END r0_rd_out[379]
  PIN r0_rd_out[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 125.199 165.870 125.217 165.888 ;
    END
  END r0_rd_out[380]
  PIN r0_rd_out[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 126.207 165.870 126.225 165.888 ;
    END
  END r0_rd_out[381]
  PIN r0_rd_out[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 127.215 165.870 127.233 165.888 ;
    END
  END r0_rd_out[382]
  PIN r0_rd_out[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 128.223 165.870 128.241 165.888 ;
    END
  END r0_rd_out[383]
  PIN r0_rd_out[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 129.231 165.870 129.249 165.888 ;
    END
  END r0_rd_out[384]
  PIN r0_rd_out[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 130.239 165.870 130.257 165.888 ;
    END
  END r0_rd_out[385]
  PIN r0_rd_out[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 131.247 165.870 131.265 165.888 ;
    END
  END r0_rd_out[386]
  PIN r0_rd_out[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 132.255 165.870 132.273 165.888 ;
    END
  END r0_rd_out[387]
  PIN r0_rd_out[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 133.263 165.870 133.281 165.888 ;
    END
  END r0_rd_out[388]
  PIN r0_rd_out[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 134.271 165.870 134.289 165.888 ;
    END
  END r0_rd_out[389]
  PIN r0_rd_out[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 135.279 165.870 135.297 165.888 ;
    END
  END r0_rd_out[390]
  PIN r0_rd_out[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 136.287 165.870 136.305 165.888 ;
    END
  END r0_rd_out[391]
  PIN r0_rd_out[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 137.295 165.870 137.313 165.888 ;
    END
  END r0_rd_out[392]
  PIN r0_rd_out[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 138.303 165.870 138.321 165.888 ;
    END
  END r0_rd_out[393]
  PIN r0_rd_out[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 139.311 165.870 139.329 165.888 ;
    END
  END r0_rd_out[394]
  PIN r0_rd_out[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 140.319 165.870 140.337 165.888 ;
    END
  END r0_rd_out[395]
  PIN r0_rd_out[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 141.327 165.870 141.345 165.888 ;
    END
  END r0_rd_out[396]
  PIN r0_rd_out[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 142.335 165.870 142.353 165.888 ;
    END
  END r0_rd_out[397]
  PIN r0_rd_out[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 143.343 165.870 143.361 165.888 ;
    END
  END r0_rd_out[398]
  PIN r0_rd_out[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 144.351 165.870 144.369 165.888 ;
    END
  END r0_rd_out[399]
  PIN r0_rd_out[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 145.359 165.870 145.377 165.888 ;
    END
  END r0_rd_out[400]
  PIN r0_rd_out[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 146.367 165.870 146.385 165.888 ;
    END
  END r0_rd_out[401]
  PIN r0_rd_out[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 147.375 165.870 147.393 165.888 ;
    END
  END r0_rd_out[402]
  PIN r0_rd_out[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 148.383 165.870 148.401 165.888 ;
    END
  END r0_rd_out[403]
  PIN r0_rd_out[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 149.391 165.870 149.409 165.888 ;
    END
  END r0_rd_out[404]
  PIN r0_rd_out[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 150.399 165.870 150.417 165.888 ;
    END
  END r0_rd_out[405]
  PIN r0_rd_out[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 151.407 165.870 151.425 165.888 ;
    END
  END r0_rd_out[406]
  PIN r0_rd_out[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 152.415 165.870 152.433 165.888 ;
    END
  END r0_rd_out[407]
  PIN r0_rd_out[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 153.423 165.870 153.441 165.888 ;
    END
  END r0_rd_out[408]
  PIN r0_rd_out[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 154.431 165.870 154.449 165.888 ;
    END
  END r0_rd_out[409]
  PIN r0_rd_out[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 155.439 165.870 155.457 165.888 ;
    END
  END r0_rd_out[410]
  PIN r0_rd_out[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 156.447 165.870 156.465 165.888 ;
    END
  END r0_rd_out[411]
  PIN r0_rd_out[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 157.455 165.870 157.473 165.888 ;
    END
  END r0_rd_out[412]
  PIN r0_rd_out[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 158.463 165.870 158.481 165.888 ;
    END
  END r0_rd_out[413]
  PIN r0_rd_out[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 159.471 165.870 159.489 165.888 ;
    END
  END r0_rd_out[414]
  PIN r0_rd_out[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 160.479 165.870 160.497 165.888 ;
    END
  END r0_rd_out[415]
  PIN r0_rd_out[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 161.487 165.870 161.505 165.888 ;
    END
  END r0_rd_out[416]
  PIN r0_rd_out[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 162.495 165.870 162.513 165.888 ;
    END
  END r0_rd_out[417]
  PIN r0_rd_out[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 163.503 165.870 163.521 165.888 ;
    END
  END r0_rd_out[418]
  PIN r0_rd_out[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 164.511 165.870 164.529 165.888 ;
    END
  END r0_rd_out[419]
  PIN r0_rd_out[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 165.519 165.870 165.537 165.888 ;
    END
  END r0_rd_out[420]
  PIN r0_rd_out[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 166.527 165.870 166.545 165.888 ;
    END
  END r0_rd_out[421]
  PIN r0_rd_out[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 167.535 165.870 167.553 165.888 ;
    END
  END r0_rd_out[422]
  PIN r0_rd_out[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 168.543 165.870 168.561 165.888 ;
    END
  END r0_rd_out[423]
  PIN r0_rd_out[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 169.551 165.870 169.569 165.888 ;
    END
  END r0_rd_out[424]
  PIN r0_rd_out[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 170.559 165.870 170.577 165.888 ;
    END
  END r0_rd_out[425]
  PIN r0_rd_out[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 171.567 165.870 171.585 165.888 ;
    END
  END r0_rd_out[426]
  PIN r0_rd_out[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 172.575 165.870 172.593 165.888 ;
    END
  END r0_rd_out[427]
  PIN r0_rd_out[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 173.583 165.870 173.601 165.888 ;
    END
  END r0_rd_out[428]
  PIN r0_rd_out[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 174.591 165.870 174.609 165.888 ;
    END
  END r0_rd_out[429]
  PIN r0_rd_out[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 175.599 165.870 175.617 165.888 ;
    END
  END r0_rd_out[430]
  PIN r0_rd_out[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 176.607 165.870 176.625 165.888 ;
    END
  END r0_rd_out[431]
  PIN r0_rd_out[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 177.615 165.870 177.633 165.888 ;
    END
  END r0_rd_out[432]
  PIN r0_rd_out[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 178.623 165.870 178.641 165.888 ;
    END
  END r0_rd_out[433]
  PIN r0_rd_out[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 179.631 165.870 179.649 165.888 ;
    END
  END r0_rd_out[434]
  PIN r0_rd_out[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 180.639 165.870 180.657 165.888 ;
    END
  END r0_rd_out[435]
  PIN r0_rd_out[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 181.647 165.870 181.665 165.888 ;
    END
  END r0_rd_out[436]
  PIN r0_rd_out[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 182.655 165.870 182.673 165.888 ;
    END
  END r0_rd_out[437]
  PIN r0_rd_out[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 183.663 165.870 183.681 165.888 ;
    END
  END r0_rd_out[438]
  PIN r0_rd_out[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 184.671 165.870 184.689 165.888 ;
    END
  END r0_rd_out[439]
  PIN r0_rd_out[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 185.679 165.870 185.697 165.888 ;
    END
  END r0_rd_out[440]
  PIN r0_rd_out[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 186.687 165.870 186.705 165.888 ;
    END
  END r0_rd_out[441]
  PIN r0_rd_out[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 187.695 165.870 187.713 165.888 ;
    END
  END r0_rd_out[442]
  PIN r0_rd_out[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 188.703 165.870 188.721 165.888 ;
    END
  END r0_rd_out[443]
  PIN r0_rd_out[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 189.711 165.870 189.729 165.888 ;
    END
  END r0_rd_out[444]
  PIN r0_rd_out[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 190.719 165.870 190.737 165.888 ;
    END
  END r0_rd_out[445]
  PIN r0_rd_out[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 191.727 165.870 191.745 165.888 ;
    END
  END r0_rd_out[446]
  PIN r0_rd_out[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 192.735 165.870 192.753 165.888 ;
    END
  END r0_rd_out[447]
  PIN r0_rd_out[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 193.743 165.870 193.761 165.888 ;
    END
  END r0_rd_out[448]
  PIN r0_rd_out[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 194.751 165.870 194.769 165.888 ;
    END
  END r0_rd_out[449]
  PIN r0_rd_out[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 195.759 165.870 195.777 165.888 ;
    END
  END r0_rd_out[450]
  PIN r0_rd_out[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 196.767 165.870 196.785 165.888 ;
    END
  END r0_rd_out[451]
  PIN r0_rd_out[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 197.775 165.870 197.793 165.888 ;
    END
  END r0_rd_out[452]
  PIN r0_rd_out[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 198.783 165.870 198.801 165.888 ;
    END
  END r0_rd_out[453]
  PIN r0_rd_out[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 199.791 165.870 199.809 165.888 ;
    END
  END r0_rd_out[454]
  PIN r0_rd_out[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 200.799 165.870 200.817 165.888 ;
    END
  END r0_rd_out[455]
  PIN r0_rd_out[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 201.807 165.870 201.825 165.888 ;
    END
  END r0_rd_out[456]
  PIN r0_rd_out[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 202.815 165.870 202.833 165.888 ;
    END
  END r0_rd_out[457]
  PIN r0_rd_out[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 203.823 165.870 203.841 165.888 ;
    END
  END r0_rd_out[458]
  PIN r0_rd_out[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 204.831 165.870 204.849 165.888 ;
    END
  END r0_rd_out[459]
  PIN r0_rd_out[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 205.839 165.870 205.857 165.888 ;
    END
  END r0_rd_out[460]
  PIN r0_rd_out[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 206.847 165.870 206.865 165.888 ;
    END
  END r0_rd_out[461]
  PIN r0_rd_out[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 207.855 165.870 207.873 165.888 ;
    END
  END r0_rd_out[462]
  PIN r0_rd_out[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 208.863 165.870 208.881 165.888 ;
    END
  END r0_rd_out[463]
  PIN r0_rd_out[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 209.871 165.870 209.889 165.888 ;
    END
  END r0_rd_out[464]
  PIN r0_rd_out[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 210.879 165.870 210.897 165.888 ;
    END
  END r0_rd_out[465]
  PIN r0_rd_out[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 211.887 165.870 211.905 165.888 ;
    END
  END r0_rd_out[466]
  PIN r0_rd_out[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 212.895 165.870 212.913 165.888 ;
    END
  END r0_rd_out[467]
  PIN r0_rd_out[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 213.903 165.870 213.921 165.888 ;
    END
  END r0_rd_out[468]
  PIN r0_rd_out[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 214.911 165.870 214.929 165.888 ;
    END
  END r0_rd_out[469]
  PIN r0_rd_out[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 215.919 165.870 215.937 165.888 ;
    END
  END r0_rd_out[470]
  PIN r0_rd_out[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 216.927 165.870 216.945 165.888 ;
    END
  END r0_rd_out[471]
  PIN r0_rd_out[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 217.935 165.870 217.953 165.888 ;
    END
  END r0_rd_out[472]
  PIN r0_rd_out[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 218.943 165.870 218.961 165.888 ;
    END
  END r0_rd_out[473]
  PIN r0_rd_out[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 219.951 165.870 219.969 165.888 ;
    END
  END r0_rd_out[474]
  PIN r0_rd_out[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 220.959 165.870 220.977 165.888 ;
    END
  END r0_rd_out[475]
  PIN r0_rd_out[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 221.967 165.870 221.985 165.888 ;
    END
  END r0_rd_out[476]
  PIN r0_rd_out[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 222.975 165.870 222.993 165.888 ;
    END
  END r0_rd_out[477]
  PIN r0_rd_out[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 223.983 165.870 224.001 165.888 ;
    END
  END r0_rd_out[478]
  PIN r0_rd_out[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 224.991 165.870 225.009 165.888 ;
    END
  END r0_rd_out[479]
  PIN r0_rd_out[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 225.999 165.870 226.017 165.888 ;
    END
  END r0_rd_out[480]
  PIN r0_rd_out[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 227.007 165.870 227.025 165.888 ;
    END
  END r0_rd_out[481]
  PIN r0_rd_out[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 228.015 165.870 228.033 165.888 ;
    END
  END r0_rd_out[482]
  PIN r0_rd_out[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 229.023 165.870 229.041 165.888 ;
    END
  END r0_rd_out[483]
  PIN r0_rd_out[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 230.031 165.870 230.049 165.888 ;
    END
  END r0_rd_out[484]
  PIN r0_rd_out[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 231.039 165.870 231.057 165.888 ;
    END
  END r0_rd_out[485]
  PIN r0_rd_out[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 232.047 165.870 232.065 165.888 ;
    END
  END r0_rd_out[486]
  PIN r0_rd_out[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 233.055 165.870 233.073 165.888 ;
    END
  END r0_rd_out[487]
  PIN r0_rd_out[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 234.063 165.870 234.081 165.888 ;
    END
  END r0_rd_out[488]
  PIN r0_rd_out[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 235.071 165.870 235.089 165.888 ;
    END
  END r0_rd_out[489]
  PIN r0_rd_out[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 236.079 165.870 236.097 165.888 ;
    END
  END r0_rd_out[490]
  PIN r0_rd_out[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 237.087 165.870 237.105 165.888 ;
    END
  END r0_rd_out[491]
  PIN r0_rd_out[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 238.095 165.870 238.113 165.888 ;
    END
  END r0_rd_out[492]
  PIN r0_rd_out[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 239.103 165.870 239.121 165.888 ;
    END
  END r0_rd_out[493]
  PIN r0_rd_out[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 240.111 165.870 240.129 165.888 ;
    END
  END r0_rd_out[494]
  PIN r0_rd_out[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 241.119 165.870 241.137 165.888 ;
    END
  END r0_rd_out[495]
  PIN r0_rd_out[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 242.127 165.870 242.145 165.888 ;
    END
  END r0_rd_out[496]
  PIN r0_rd_out[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 243.135 165.870 243.153 165.888 ;
    END
  END r0_rd_out[497]
  PIN r0_rd_out[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 244.143 165.870 244.161 165.888 ;
    END
  END r0_rd_out[498]
  PIN r0_rd_out[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 245.151 165.870 245.169 165.888 ;
    END
  END r0_rd_out[499]
  PIN r0_rd_out[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 246.159 165.870 246.177 165.888 ;
    END
  END r0_rd_out[500]
  PIN r0_rd_out[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 247.167 165.870 247.185 165.888 ;
    END
  END r0_rd_out[501]
  PIN r0_rd_out[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 248.175 165.870 248.193 165.888 ;
    END
  END r0_rd_out[502]
  PIN r0_rd_out[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 249.183 165.870 249.201 165.888 ;
    END
  END r0_rd_out[503]
  PIN r0_rd_out[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 250.191 165.870 250.209 165.888 ;
    END
  END r0_rd_out[504]
  PIN r0_rd_out[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 251.199 165.870 251.217 165.888 ;
    END
  END r0_rd_out[505]
  PIN r0_rd_out[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 252.207 165.870 252.225 165.888 ;
    END
  END r0_rd_out[506]
  PIN r0_rd_out[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 253.215 165.870 253.233 165.888 ;
    END
  END r0_rd_out[507]
  PIN r0_rd_out[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 254.223 165.870 254.241 165.888 ;
    END
  END r0_rd_out[508]
  PIN r0_rd_out[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 255.231 165.870 255.249 165.888 ;
    END
  END r0_rd_out[509]
  PIN r0_rd_out[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 256.239 165.870 256.257 165.888 ;
    END
  END r0_rd_out[510]
  PIN r0_rd_out[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 257.247 165.870 257.265 165.888 ;
    END
  END r0_rd_out[511]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 147.732 0.024 147.756 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 148.884 0.024 148.908 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 150.036 0.024 150.060 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 151.188 0.024 151.212 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 152.340 0.024 152.364 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 153.492 0.024 153.516 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 147.732 265.421 147.756 ;
    END
  END w0_addr_in[6]
  PIN w0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 148.884 265.421 148.908 ;
    END
  END w0_addr_in[7]
  PIN w0_addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 150.036 265.421 150.060 ;
    END
  END w0_addr_in[8]
  PIN w0_addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 151.188 265.421 151.212 ;
    END
  END w0_addr_in[9]
  PIN w0_addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 152.340 265.421 152.364 ;
    END
  END w0_addr_in[10]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 154.644 0.024 154.668 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 155.796 0.024 155.820 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 156.948 0.024 156.972 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 158.100 0.024 158.124 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 159.252 0.024 159.276 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 160.404 0.024 160.428 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 153.492 265.421 153.516 ;
    END
  END r0_addr_in[6]
  PIN r0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 154.644 265.421 154.668 ;
    END
  END r0_addr_in[7]
  PIN r0_addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 155.796 265.421 155.820 ;
    END
  END r0_addr_in[8]
  PIN r0_addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 156.948 265.421 156.972 ;
    END
  END r0_addr_in[9]
  PIN r0_addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.397 158.100 265.421 158.124 ;
    END
  END r0_addr_in[10]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 258.255 165.870 258.273 165.888 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 259.263 165.870 259.281 165.888 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 260.271 165.870 260.289 165.888 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 261.279 165.870 261.297 165.888 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 262.287 165.870 262.305 165.888 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.108 0.192 265.313 0.288 ;
      RECT 0.108 0.960 265.313 1.056 ;
      RECT 0.108 1.728 265.313 1.824 ;
      RECT 0.108 2.496 265.313 2.592 ;
      RECT 0.108 3.264 265.313 3.360 ;
      RECT 0.108 4.032 265.313 4.128 ;
      RECT 0.108 4.800 265.313 4.896 ;
      RECT 0.108 5.568 265.313 5.664 ;
      RECT 0.108 6.336 265.313 6.432 ;
      RECT 0.108 7.104 265.313 7.200 ;
      RECT 0.108 7.872 265.313 7.968 ;
      RECT 0.108 8.640 265.313 8.736 ;
      RECT 0.108 9.408 265.313 9.504 ;
      RECT 0.108 10.176 265.313 10.272 ;
      RECT 0.108 10.944 265.313 11.040 ;
      RECT 0.108 11.712 265.313 11.808 ;
      RECT 0.108 12.480 265.313 12.576 ;
      RECT 0.108 13.248 265.313 13.344 ;
      RECT 0.108 14.016 265.313 14.112 ;
      RECT 0.108 14.784 265.313 14.880 ;
      RECT 0.108 15.552 265.313 15.648 ;
      RECT 0.108 16.320 265.313 16.416 ;
      RECT 0.108 17.088 265.313 17.184 ;
      RECT 0.108 17.856 265.313 17.952 ;
      RECT 0.108 18.624 265.313 18.720 ;
      RECT 0.108 19.392 265.313 19.488 ;
      RECT 0.108 20.160 265.313 20.256 ;
      RECT 0.108 20.928 265.313 21.024 ;
      RECT 0.108 21.696 265.313 21.792 ;
      RECT 0.108 22.464 265.313 22.560 ;
      RECT 0.108 23.232 265.313 23.328 ;
      RECT 0.108 24.000 265.313 24.096 ;
      RECT 0.108 24.768 265.313 24.864 ;
      RECT 0.108 25.536 265.313 25.632 ;
      RECT 0.108 26.304 265.313 26.400 ;
      RECT 0.108 27.072 265.313 27.168 ;
      RECT 0.108 27.840 265.313 27.936 ;
      RECT 0.108 28.608 265.313 28.704 ;
      RECT 0.108 29.376 265.313 29.472 ;
      RECT 0.108 30.144 265.313 30.240 ;
      RECT 0.108 30.912 265.313 31.008 ;
      RECT 0.108 31.680 265.313 31.776 ;
      RECT 0.108 32.448 265.313 32.544 ;
      RECT 0.108 33.216 265.313 33.312 ;
      RECT 0.108 33.984 265.313 34.080 ;
      RECT 0.108 34.752 265.313 34.848 ;
      RECT 0.108 35.520 265.313 35.616 ;
      RECT 0.108 36.288 265.313 36.384 ;
      RECT 0.108 37.056 265.313 37.152 ;
      RECT 0.108 37.824 265.313 37.920 ;
      RECT 0.108 38.592 265.313 38.688 ;
      RECT 0.108 39.360 265.313 39.456 ;
      RECT 0.108 40.128 265.313 40.224 ;
      RECT 0.108 40.896 265.313 40.992 ;
      RECT 0.108 41.664 265.313 41.760 ;
      RECT 0.108 42.432 265.313 42.528 ;
      RECT 0.108 43.200 265.313 43.296 ;
      RECT 0.108 43.968 265.313 44.064 ;
      RECT 0.108 44.736 265.313 44.832 ;
      RECT 0.108 45.504 265.313 45.600 ;
      RECT 0.108 46.272 265.313 46.368 ;
      RECT 0.108 47.040 265.313 47.136 ;
      RECT 0.108 47.808 265.313 47.904 ;
      RECT 0.108 48.576 265.313 48.672 ;
      RECT 0.108 49.344 265.313 49.440 ;
      RECT 0.108 50.112 265.313 50.208 ;
      RECT 0.108 50.880 265.313 50.976 ;
      RECT 0.108 51.648 265.313 51.744 ;
      RECT 0.108 52.416 265.313 52.512 ;
      RECT 0.108 53.184 265.313 53.280 ;
      RECT 0.108 53.952 265.313 54.048 ;
      RECT 0.108 54.720 265.313 54.816 ;
      RECT 0.108 55.488 265.313 55.584 ;
      RECT 0.108 56.256 265.313 56.352 ;
      RECT 0.108 57.024 265.313 57.120 ;
      RECT 0.108 57.792 265.313 57.888 ;
      RECT 0.108 58.560 265.313 58.656 ;
      RECT 0.108 59.328 265.313 59.424 ;
      RECT 0.108 60.096 265.313 60.192 ;
      RECT 0.108 60.864 265.313 60.960 ;
      RECT 0.108 61.632 265.313 61.728 ;
      RECT 0.108 62.400 265.313 62.496 ;
      RECT 0.108 63.168 265.313 63.264 ;
      RECT 0.108 63.936 265.313 64.032 ;
      RECT 0.108 64.704 265.313 64.800 ;
      RECT 0.108 65.472 265.313 65.568 ;
      RECT 0.108 66.240 265.313 66.336 ;
      RECT 0.108 67.008 265.313 67.104 ;
      RECT 0.108 67.776 265.313 67.872 ;
      RECT 0.108 68.544 265.313 68.640 ;
      RECT 0.108 69.312 265.313 69.408 ;
      RECT 0.108 70.080 265.313 70.176 ;
      RECT 0.108 70.848 265.313 70.944 ;
      RECT 0.108 71.616 265.313 71.712 ;
      RECT 0.108 72.384 265.313 72.480 ;
      RECT 0.108 73.152 265.313 73.248 ;
      RECT 0.108 73.920 265.313 74.016 ;
      RECT 0.108 74.688 265.313 74.784 ;
      RECT 0.108 75.456 265.313 75.552 ;
      RECT 0.108 76.224 265.313 76.320 ;
      RECT 0.108 76.992 265.313 77.088 ;
      RECT 0.108 77.760 265.313 77.856 ;
      RECT 0.108 78.528 265.313 78.624 ;
      RECT 0.108 79.296 265.313 79.392 ;
      RECT 0.108 80.064 265.313 80.160 ;
      RECT 0.108 80.832 265.313 80.928 ;
      RECT 0.108 81.600 265.313 81.696 ;
      RECT 0.108 82.368 265.313 82.464 ;
      RECT 0.108 83.136 265.313 83.232 ;
      RECT 0.108 83.904 265.313 84.000 ;
      RECT 0.108 84.672 265.313 84.768 ;
      RECT 0.108 85.440 265.313 85.536 ;
      RECT 0.108 86.208 265.313 86.304 ;
      RECT 0.108 86.976 265.313 87.072 ;
      RECT 0.108 87.744 265.313 87.840 ;
      RECT 0.108 88.512 265.313 88.608 ;
      RECT 0.108 89.280 265.313 89.376 ;
      RECT 0.108 90.048 265.313 90.144 ;
      RECT 0.108 90.816 265.313 90.912 ;
      RECT 0.108 91.584 265.313 91.680 ;
      RECT 0.108 92.352 265.313 92.448 ;
      RECT 0.108 93.120 265.313 93.216 ;
      RECT 0.108 93.888 265.313 93.984 ;
      RECT 0.108 94.656 265.313 94.752 ;
      RECT 0.108 95.424 265.313 95.520 ;
      RECT 0.108 96.192 265.313 96.288 ;
      RECT 0.108 96.960 265.313 97.056 ;
      RECT 0.108 97.728 265.313 97.824 ;
      RECT 0.108 98.496 265.313 98.592 ;
      RECT 0.108 99.264 265.313 99.360 ;
      RECT 0.108 100.032 265.313 100.128 ;
      RECT 0.108 100.800 265.313 100.896 ;
      RECT 0.108 101.568 265.313 101.664 ;
      RECT 0.108 102.336 265.313 102.432 ;
      RECT 0.108 103.104 265.313 103.200 ;
      RECT 0.108 103.872 265.313 103.968 ;
      RECT 0.108 104.640 265.313 104.736 ;
      RECT 0.108 105.408 265.313 105.504 ;
      RECT 0.108 106.176 265.313 106.272 ;
      RECT 0.108 106.944 265.313 107.040 ;
      RECT 0.108 107.712 265.313 107.808 ;
      RECT 0.108 108.480 265.313 108.576 ;
      RECT 0.108 109.248 265.313 109.344 ;
      RECT 0.108 110.016 265.313 110.112 ;
      RECT 0.108 110.784 265.313 110.880 ;
      RECT 0.108 111.552 265.313 111.648 ;
      RECT 0.108 112.320 265.313 112.416 ;
      RECT 0.108 113.088 265.313 113.184 ;
      RECT 0.108 113.856 265.313 113.952 ;
      RECT 0.108 114.624 265.313 114.720 ;
      RECT 0.108 115.392 265.313 115.488 ;
      RECT 0.108 116.160 265.313 116.256 ;
      RECT 0.108 116.928 265.313 117.024 ;
      RECT 0.108 117.696 265.313 117.792 ;
      RECT 0.108 118.464 265.313 118.560 ;
      RECT 0.108 119.232 265.313 119.328 ;
      RECT 0.108 120.000 265.313 120.096 ;
      RECT 0.108 120.768 265.313 120.864 ;
      RECT 0.108 121.536 265.313 121.632 ;
      RECT 0.108 122.304 265.313 122.400 ;
      RECT 0.108 123.072 265.313 123.168 ;
      RECT 0.108 123.840 265.313 123.936 ;
      RECT 0.108 124.608 265.313 124.704 ;
      RECT 0.108 125.376 265.313 125.472 ;
      RECT 0.108 126.144 265.313 126.240 ;
      RECT 0.108 126.912 265.313 127.008 ;
      RECT 0.108 127.680 265.313 127.776 ;
      RECT 0.108 128.448 265.313 128.544 ;
      RECT 0.108 129.216 265.313 129.312 ;
      RECT 0.108 129.984 265.313 130.080 ;
      RECT 0.108 130.752 265.313 130.848 ;
      RECT 0.108 131.520 265.313 131.616 ;
      RECT 0.108 132.288 265.313 132.384 ;
      RECT 0.108 133.056 265.313 133.152 ;
      RECT 0.108 133.824 265.313 133.920 ;
      RECT 0.108 134.592 265.313 134.688 ;
      RECT 0.108 135.360 265.313 135.456 ;
      RECT 0.108 136.128 265.313 136.224 ;
      RECT 0.108 136.896 265.313 136.992 ;
      RECT 0.108 137.664 265.313 137.760 ;
      RECT 0.108 138.432 265.313 138.528 ;
      RECT 0.108 139.200 265.313 139.296 ;
      RECT 0.108 139.968 265.313 140.064 ;
      RECT 0.108 140.736 265.313 140.832 ;
      RECT 0.108 141.504 265.313 141.600 ;
      RECT 0.108 142.272 265.313 142.368 ;
      RECT 0.108 143.040 265.313 143.136 ;
      RECT 0.108 143.808 265.313 143.904 ;
      RECT 0.108 144.576 265.313 144.672 ;
      RECT 0.108 145.344 265.313 145.440 ;
      RECT 0.108 146.112 265.313 146.208 ;
      RECT 0.108 146.880 265.313 146.976 ;
      RECT 0.108 147.648 265.313 147.744 ;
      RECT 0.108 148.416 265.313 148.512 ;
      RECT 0.108 149.184 265.313 149.280 ;
      RECT 0.108 149.952 265.313 150.048 ;
      RECT 0.108 150.720 265.313 150.816 ;
      RECT 0.108 151.488 265.313 151.584 ;
      RECT 0.108 152.256 265.313 152.352 ;
      RECT 0.108 153.024 265.313 153.120 ;
      RECT 0.108 153.792 265.313 153.888 ;
      RECT 0.108 154.560 265.313 154.656 ;
      RECT 0.108 155.328 265.313 155.424 ;
      RECT 0.108 156.096 265.313 156.192 ;
      RECT 0.108 156.864 265.313 156.960 ;
      RECT 0.108 157.632 265.313 157.728 ;
      RECT 0.108 158.400 265.313 158.496 ;
      RECT 0.108 159.168 265.313 159.264 ;
      RECT 0.108 159.936 265.313 160.032 ;
      RECT 0.108 160.704 265.313 160.800 ;
      RECT 0.108 161.472 265.313 161.568 ;
      RECT 0.108 162.240 265.313 162.336 ;
      RECT 0.108 163.008 265.313 163.104 ;
      RECT 0.108 163.776 265.313 163.872 ;
      RECT 0.108 164.544 265.313 164.640 ;
      RECT 0.108 165.312 265.313 165.408 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.108 0.192 265.313 0.288 ;
      RECT 0.108 0.960 265.313 1.056 ;
      RECT 0.108 1.728 265.313 1.824 ;
      RECT 0.108 2.496 265.313 2.592 ;
      RECT 0.108 3.264 265.313 3.360 ;
      RECT 0.108 4.032 265.313 4.128 ;
      RECT 0.108 4.800 265.313 4.896 ;
      RECT 0.108 5.568 265.313 5.664 ;
      RECT 0.108 6.336 265.313 6.432 ;
      RECT 0.108 7.104 265.313 7.200 ;
      RECT 0.108 7.872 265.313 7.968 ;
      RECT 0.108 8.640 265.313 8.736 ;
      RECT 0.108 9.408 265.313 9.504 ;
      RECT 0.108 10.176 265.313 10.272 ;
      RECT 0.108 10.944 265.313 11.040 ;
      RECT 0.108 11.712 265.313 11.808 ;
      RECT 0.108 12.480 265.313 12.576 ;
      RECT 0.108 13.248 265.313 13.344 ;
      RECT 0.108 14.016 265.313 14.112 ;
      RECT 0.108 14.784 265.313 14.880 ;
      RECT 0.108 15.552 265.313 15.648 ;
      RECT 0.108 16.320 265.313 16.416 ;
      RECT 0.108 17.088 265.313 17.184 ;
      RECT 0.108 17.856 265.313 17.952 ;
      RECT 0.108 18.624 265.313 18.720 ;
      RECT 0.108 19.392 265.313 19.488 ;
      RECT 0.108 20.160 265.313 20.256 ;
      RECT 0.108 20.928 265.313 21.024 ;
      RECT 0.108 21.696 265.313 21.792 ;
      RECT 0.108 22.464 265.313 22.560 ;
      RECT 0.108 23.232 265.313 23.328 ;
      RECT 0.108 24.000 265.313 24.096 ;
      RECT 0.108 24.768 265.313 24.864 ;
      RECT 0.108 25.536 265.313 25.632 ;
      RECT 0.108 26.304 265.313 26.400 ;
      RECT 0.108 27.072 265.313 27.168 ;
      RECT 0.108 27.840 265.313 27.936 ;
      RECT 0.108 28.608 265.313 28.704 ;
      RECT 0.108 29.376 265.313 29.472 ;
      RECT 0.108 30.144 265.313 30.240 ;
      RECT 0.108 30.912 265.313 31.008 ;
      RECT 0.108 31.680 265.313 31.776 ;
      RECT 0.108 32.448 265.313 32.544 ;
      RECT 0.108 33.216 265.313 33.312 ;
      RECT 0.108 33.984 265.313 34.080 ;
      RECT 0.108 34.752 265.313 34.848 ;
      RECT 0.108 35.520 265.313 35.616 ;
      RECT 0.108 36.288 265.313 36.384 ;
      RECT 0.108 37.056 265.313 37.152 ;
      RECT 0.108 37.824 265.313 37.920 ;
      RECT 0.108 38.592 265.313 38.688 ;
      RECT 0.108 39.360 265.313 39.456 ;
      RECT 0.108 40.128 265.313 40.224 ;
      RECT 0.108 40.896 265.313 40.992 ;
      RECT 0.108 41.664 265.313 41.760 ;
      RECT 0.108 42.432 265.313 42.528 ;
      RECT 0.108 43.200 265.313 43.296 ;
      RECT 0.108 43.968 265.313 44.064 ;
      RECT 0.108 44.736 265.313 44.832 ;
      RECT 0.108 45.504 265.313 45.600 ;
      RECT 0.108 46.272 265.313 46.368 ;
      RECT 0.108 47.040 265.313 47.136 ;
      RECT 0.108 47.808 265.313 47.904 ;
      RECT 0.108 48.576 265.313 48.672 ;
      RECT 0.108 49.344 265.313 49.440 ;
      RECT 0.108 50.112 265.313 50.208 ;
      RECT 0.108 50.880 265.313 50.976 ;
      RECT 0.108 51.648 265.313 51.744 ;
      RECT 0.108 52.416 265.313 52.512 ;
      RECT 0.108 53.184 265.313 53.280 ;
      RECT 0.108 53.952 265.313 54.048 ;
      RECT 0.108 54.720 265.313 54.816 ;
      RECT 0.108 55.488 265.313 55.584 ;
      RECT 0.108 56.256 265.313 56.352 ;
      RECT 0.108 57.024 265.313 57.120 ;
      RECT 0.108 57.792 265.313 57.888 ;
      RECT 0.108 58.560 265.313 58.656 ;
      RECT 0.108 59.328 265.313 59.424 ;
      RECT 0.108 60.096 265.313 60.192 ;
      RECT 0.108 60.864 265.313 60.960 ;
      RECT 0.108 61.632 265.313 61.728 ;
      RECT 0.108 62.400 265.313 62.496 ;
      RECT 0.108 63.168 265.313 63.264 ;
      RECT 0.108 63.936 265.313 64.032 ;
      RECT 0.108 64.704 265.313 64.800 ;
      RECT 0.108 65.472 265.313 65.568 ;
      RECT 0.108 66.240 265.313 66.336 ;
      RECT 0.108 67.008 265.313 67.104 ;
      RECT 0.108 67.776 265.313 67.872 ;
      RECT 0.108 68.544 265.313 68.640 ;
      RECT 0.108 69.312 265.313 69.408 ;
      RECT 0.108 70.080 265.313 70.176 ;
      RECT 0.108 70.848 265.313 70.944 ;
      RECT 0.108 71.616 265.313 71.712 ;
      RECT 0.108 72.384 265.313 72.480 ;
      RECT 0.108 73.152 265.313 73.248 ;
      RECT 0.108 73.920 265.313 74.016 ;
      RECT 0.108 74.688 265.313 74.784 ;
      RECT 0.108 75.456 265.313 75.552 ;
      RECT 0.108 76.224 265.313 76.320 ;
      RECT 0.108 76.992 265.313 77.088 ;
      RECT 0.108 77.760 265.313 77.856 ;
      RECT 0.108 78.528 265.313 78.624 ;
      RECT 0.108 79.296 265.313 79.392 ;
      RECT 0.108 80.064 265.313 80.160 ;
      RECT 0.108 80.832 265.313 80.928 ;
      RECT 0.108 81.600 265.313 81.696 ;
      RECT 0.108 82.368 265.313 82.464 ;
      RECT 0.108 83.136 265.313 83.232 ;
      RECT 0.108 83.904 265.313 84.000 ;
      RECT 0.108 84.672 265.313 84.768 ;
      RECT 0.108 85.440 265.313 85.536 ;
      RECT 0.108 86.208 265.313 86.304 ;
      RECT 0.108 86.976 265.313 87.072 ;
      RECT 0.108 87.744 265.313 87.840 ;
      RECT 0.108 88.512 265.313 88.608 ;
      RECT 0.108 89.280 265.313 89.376 ;
      RECT 0.108 90.048 265.313 90.144 ;
      RECT 0.108 90.816 265.313 90.912 ;
      RECT 0.108 91.584 265.313 91.680 ;
      RECT 0.108 92.352 265.313 92.448 ;
      RECT 0.108 93.120 265.313 93.216 ;
      RECT 0.108 93.888 265.313 93.984 ;
      RECT 0.108 94.656 265.313 94.752 ;
      RECT 0.108 95.424 265.313 95.520 ;
      RECT 0.108 96.192 265.313 96.288 ;
      RECT 0.108 96.960 265.313 97.056 ;
      RECT 0.108 97.728 265.313 97.824 ;
      RECT 0.108 98.496 265.313 98.592 ;
      RECT 0.108 99.264 265.313 99.360 ;
      RECT 0.108 100.032 265.313 100.128 ;
      RECT 0.108 100.800 265.313 100.896 ;
      RECT 0.108 101.568 265.313 101.664 ;
      RECT 0.108 102.336 265.313 102.432 ;
      RECT 0.108 103.104 265.313 103.200 ;
      RECT 0.108 103.872 265.313 103.968 ;
      RECT 0.108 104.640 265.313 104.736 ;
      RECT 0.108 105.408 265.313 105.504 ;
      RECT 0.108 106.176 265.313 106.272 ;
      RECT 0.108 106.944 265.313 107.040 ;
      RECT 0.108 107.712 265.313 107.808 ;
      RECT 0.108 108.480 265.313 108.576 ;
      RECT 0.108 109.248 265.313 109.344 ;
      RECT 0.108 110.016 265.313 110.112 ;
      RECT 0.108 110.784 265.313 110.880 ;
      RECT 0.108 111.552 265.313 111.648 ;
      RECT 0.108 112.320 265.313 112.416 ;
      RECT 0.108 113.088 265.313 113.184 ;
      RECT 0.108 113.856 265.313 113.952 ;
      RECT 0.108 114.624 265.313 114.720 ;
      RECT 0.108 115.392 265.313 115.488 ;
      RECT 0.108 116.160 265.313 116.256 ;
      RECT 0.108 116.928 265.313 117.024 ;
      RECT 0.108 117.696 265.313 117.792 ;
      RECT 0.108 118.464 265.313 118.560 ;
      RECT 0.108 119.232 265.313 119.328 ;
      RECT 0.108 120.000 265.313 120.096 ;
      RECT 0.108 120.768 265.313 120.864 ;
      RECT 0.108 121.536 265.313 121.632 ;
      RECT 0.108 122.304 265.313 122.400 ;
      RECT 0.108 123.072 265.313 123.168 ;
      RECT 0.108 123.840 265.313 123.936 ;
      RECT 0.108 124.608 265.313 124.704 ;
      RECT 0.108 125.376 265.313 125.472 ;
      RECT 0.108 126.144 265.313 126.240 ;
      RECT 0.108 126.912 265.313 127.008 ;
      RECT 0.108 127.680 265.313 127.776 ;
      RECT 0.108 128.448 265.313 128.544 ;
      RECT 0.108 129.216 265.313 129.312 ;
      RECT 0.108 129.984 265.313 130.080 ;
      RECT 0.108 130.752 265.313 130.848 ;
      RECT 0.108 131.520 265.313 131.616 ;
      RECT 0.108 132.288 265.313 132.384 ;
      RECT 0.108 133.056 265.313 133.152 ;
      RECT 0.108 133.824 265.313 133.920 ;
      RECT 0.108 134.592 265.313 134.688 ;
      RECT 0.108 135.360 265.313 135.456 ;
      RECT 0.108 136.128 265.313 136.224 ;
      RECT 0.108 136.896 265.313 136.992 ;
      RECT 0.108 137.664 265.313 137.760 ;
      RECT 0.108 138.432 265.313 138.528 ;
      RECT 0.108 139.200 265.313 139.296 ;
      RECT 0.108 139.968 265.313 140.064 ;
      RECT 0.108 140.736 265.313 140.832 ;
      RECT 0.108 141.504 265.313 141.600 ;
      RECT 0.108 142.272 265.313 142.368 ;
      RECT 0.108 143.040 265.313 143.136 ;
      RECT 0.108 143.808 265.313 143.904 ;
      RECT 0.108 144.576 265.313 144.672 ;
      RECT 0.108 145.344 265.313 145.440 ;
      RECT 0.108 146.112 265.313 146.208 ;
      RECT 0.108 146.880 265.313 146.976 ;
      RECT 0.108 147.648 265.313 147.744 ;
      RECT 0.108 148.416 265.313 148.512 ;
      RECT 0.108 149.184 265.313 149.280 ;
      RECT 0.108 149.952 265.313 150.048 ;
      RECT 0.108 150.720 265.313 150.816 ;
      RECT 0.108 151.488 265.313 151.584 ;
      RECT 0.108 152.256 265.313 152.352 ;
      RECT 0.108 153.024 265.313 153.120 ;
      RECT 0.108 153.792 265.313 153.888 ;
      RECT 0.108 154.560 265.313 154.656 ;
      RECT 0.108 155.328 265.313 155.424 ;
      RECT 0.108 156.096 265.313 156.192 ;
      RECT 0.108 156.864 265.313 156.960 ;
      RECT 0.108 157.632 265.313 157.728 ;
      RECT 0.108 158.400 265.313 158.496 ;
      RECT 0.108 159.168 265.313 159.264 ;
      RECT 0.108 159.936 265.313 160.032 ;
      RECT 0.108 160.704 265.313 160.800 ;
      RECT 0.108 161.472 265.313 161.568 ;
      RECT 0.108 162.240 265.313 162.336 ;
      RECT 0.108 163.008 265.313 163.104 ;
      RECT 0.108 163.776 265.313 163.872 ;
      RECT 0.108 164.544 265.313 164.640 ;
      RECT 0.108 165.312 265.313 165.408 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 265.421 165.888 ;
    LAYER M2 ;
    RECT 0 0 265.421 165.888 ;
    LAYER M3 ;
    RECT 0 0 265.421 165.888 ;
    LAYER M4 ;
    RECT 0 0 265.421 165.888 ;
  END
END fakeram_512x2048_1r1w

END LIBRARY
