VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO liteeth_1rw1r_32w384d_8_sram
  FOREIGN liteeth_1rw1r_32w384d_8_sram 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 114.000 BY 256.200 ;
  CLASS BLOCK ;
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END clk0
  PIN csb0
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END csb0
  PIN web0
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END web0
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.045 0.070 17.115 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.925 0.070 22.995 ;
    END
  END addr0[8]
  PIN din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END din0[0]
  PIN din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END din0[1]
  PIN din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.805 0.070 28.875 ;
    END
  END din0[2]
  PIN din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.685 0.070 34.755 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END din0[9]
  PIN din0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.445 0.070 46.515 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.325 0.070 52.395 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.285 0.070 54.355 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.205 0.070 58.275 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END din0[19]
  PIN din0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.085 0.070 64.155 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.045 0.070 66.115 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.965 0.070 70.035 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.925 0.070 71.995 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.845 0.070 75.915 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.725 0.070 81.795 ;
    END
  END din0[29]
  PIN din0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.685 0.070 83.755 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END din0[31]
  PIN wmask0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.605 0.070 87.675 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.565 0.070 89.635 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.485 0.070 93.555 ;
    END
  END wmask0[3]
  PIN dout0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.445 0.070 95.515 ;
    END
  END dout0[0]
  PIN dout0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END dout0[1]
  PIN dout0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.365 0.070 99.435 ;
    END
  END dout0[2]
  PIN dout0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.325 0.070 101.395 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.285 0.070 103.355 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.245 0.070 105.315 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.205 0.070 107.275 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.125 0.070 111.195 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.085 0.070 113.155 ;
    END
  END dout0[9]
  PIN dout0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.045 0.070 115.115 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.005 0.070 117.075 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.965 0.070 119.035 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.925 0.070 120.995 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.885 0.070 122.955 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.845 0.070 124.915 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.805 0.070 126.875 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.765 0.070 128.835 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.725 0.070 130.795 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.685 0.070 132.755 ;
    END
  END dout0[19]
  PIN dout0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.645 0.070 134.715 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.605 0.070 136.675 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.565 0.070 138.635 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.525 0.070 140.595 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.485 0.070 142.555 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.445 0.070 144.515 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.405 0.070 146.475 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.365 0.070 148.435 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.325 0.070 150.395 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.285 0.070 152.355 ;
    END
  END dout0[29]
  PIN dout0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.245 0.070 154.315 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.205 0.070 156.275 ;
    END
  END dout0[31]
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.165 0.070 158.235 ;
    END
  END clk1
  PIN csb1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.125 0.070 160.195 ;
    END
  END csb1
  PIN addr1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.085 0.070 162.155 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.045 0.070 164.115 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.005 0.070 166.075 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.965 0.070 168.035 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.925 0.070 169.995 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.885 0.070 171.955 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.845 0.070 173.915 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.805 0.070 175.875 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.765 0.070 177.835 ;
    END
  END addr1[8]
  PIN dout1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.725 0.070 179.795 ;
    END
  END dout1[0]
  PIN dout1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.685 0.070 181.755 ;
    END
  END dout1[1]
  PIN dout1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.645 0.070 183.715 ;
    END
  END dout1[2]
  PIN dout1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.605 0.070 185.675 ;
    END
  END dout1[3]
  PIN dout1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.565 0.070 187.635 ;
    END
  END dout1[4]
  PIN dout1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.525 0.070 189.595 ;
    END
  END dout1[5]
  PIN dout1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.485 0.070 191.555 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.445 0.070 193.515 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.405 0.070 195.475 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.365 0.070 197.435 ;
    END
  END dout1[9]
  PIN dout1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.325 0.070 199.395 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.285 0.070 201.355 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.245 0.070 203.315 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.205 0.070 205.275 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.165 0.070 207.235 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.125 0.070 209.195 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.085 0.070 211.155 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.045 0.070 213.115 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.005 0.070 215.075 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.965 0.070 217.035 ;
    END
  END dout1[19]
  PIN dout1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.925 0.070 218.995 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.885 0.070 220.955 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.845 0.070 222.915 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.805 0.070 224.875 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.765 0.070 226.835 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.725 0.070 228.795 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.685 0.070 230.755 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.645 0.070 232.715 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.605 0.070 234.675 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.565 0.070 236.635 ;
    END
  END dout1[29]
  PIN dout1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.525 0.070 238.595 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.485 0.070 240.555 ;
    END
  END dout1[31]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 254.800 ;
      RECT 3.500 1.400 3.780 254.800 ;
      RECT 5.740 1.400 6.020 254.800 ;
      RECT 7.980 1.400 8.260 254.800 ;
      RECT 10.220 1.400 10.500 254.800 ;
      RECT 12.460 1.400 12.740 254.800 ;
      RECT 14.700 1.400 14.980 254.800 ;
      RECT 16.940 1.400 17.220 254.800 ;
      RECT 19.180 1.400 19.460 254.800 ;
      RECT 21.420 1.400 21.700 254.800 ;
      RECT 23.660 1.400 23.940 254.800 ;
      RECT 25.900 1.400 26.180 254.800 ;
      RECT 28.140 1.400 28.420 254.800 ;
      RECT 30.380 1.400 30.660 254.800 ;
      RECT 32.620 1.400 32.900 254.800 ;
      RECT 34.860 1.400 35.140 254.800 ;
      RECT 37.100 1.400 37.380 254.800 ;
      RECT 39.340 1.400 39.620 254.800 ;
      RECT 41.580 1.400 41.860 254.800 ;
      RECT 43.820 1.400 44.100 254.800 ;
      RECT 46.060 1.400 46.340 254.800 ;
      RECT 48.300 1.400 48.580 254.800 ;
      RECT 50.540 1.400 50.820 254.800 ;
      RECT 52.780 1.400 53.060 254.800 ;
      RECT 55.020 1.400 55.300 254.800 ;
      RECT 57.260 1.400 57.540 254.800 ;
      RECT 59.500 1.400 59.780 254.800 ;
      RECT 61.740 1.400 62.020 254.800 ;
      RECT 63.980 1.400 64.260 254.800 ;
      RECT 66.220 1.400 66.500 254.800 ;
      RECT 68.460 1.400 68.740 254.800 ;
      RECT 70.700 1.400 70.980 254.800 ;
      RECT 72.940 1.400 73.220 254.800 ;
      RECT 75.180 1.400 75.460 254.800 ;
      RECT 77.420 1.400 77.700 254.800 ;
      RECT 79.660 1.400 79.940 254.800 ;
      RECT 81.900 1.400 82.180 254.800 ;
      RECT 84.140 1.400 84.420 254.800 ;
      RECT 86.380 1.400 86.660 254.800 ;
      RECT 88.620 1.400 88.900 254.800 ;
      RECT 90.860 1.400 91.140 254.800 ;
      RECT 93.100 1.400 93.380 254.800 ;
      RECT 95.340 1.400 95.620 254.800 ;
      RECT 97.580 1.400 97.860 254.800 ;
      RECT 99.820 1.400 100.100 254.800 ;
      RECT 102.060 1.400 102.340 254.800 ;
      RECT 104.300 1.400 104.580 254.800 ;
      RECT 106.540 1.400 106.820 254.800 ;
      RECT 108.780 1.400 109.060 254.800 ;
      RECT 111.020 1.400 111.300 254.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 254.800 ;
      RECT 4.620 1.400 4.900 254.800 ;
      RECT 6.860 1.400 7.140 254.800 ;
      RECT 9.100 1.400 9.380 254.800 ;
      RECT 11.340 1.400 11.620 254.800 ;
      RECT 13.580 1.400 13.860 254.800 ;
      RECT 15.820 1.400 16.100 254.800 ;
      RECT 18.060 1.400 18.340 254.800 ;
      RECT 20.300 1.400 20.580 254.800 ;
      RECT 22.540 1.400 22.820 254.800 ;
      RECT 24.780 1.400 25.060 254.800 ;
      RECT 27.020 1.400 27.300 254.800 ;
      RECT 29.260 1.400 29.540 254.800 ;
      RECT 31.500 1.400 31.780 254.800 ;
      RECT 33.740 1.400 34.020 254.800 ;
      RECT 35.980 1.400 36.260 254.800 ;
      RECT 38.220 1.400 38.500 254.800 ;
      RECT 40.460 1.400 40.740 254.800 ;
      RECT 42.700 1.400 42.980 254.800 ;
      RECT 44.940 1.400 45.220 254.800 ;
      RECT 47.180 1.400 47.460 254.800 ;
      RECT 49.420 1.400 49.700 254.800 ;
      RECT 51.660 1.400 51.940 254.800 ;
      RECT 53.900 1.400 54.180 254.800 ;
      RECT 56.140 1.400 56.420 254.800 ;
      RECT 58.380 1.400 58.660 254.800 ;
      RECT 60.620 1.400 60.900 254.800 ;
      RECT 62.860 1.400 63.140 254.800 ;
      RECT 65.100 1.400 65.380 254.800 ;
      RECT 67.340 1.400 67.620 254.800 ;
      RECT 69.580 1.400 69.860 254.800 ;
      RECT 71.820 1.400 72.100 254.800 ;
      RECT 74.060 1.400 74.340 254.800 ;
      RECT 76.300 1.400 76.580 254.800 ;
      RECT 78.540 1.400 78.820 254.800 ;
      RECT 80.780 1.400 81.060 254.800 ;
      RECT 83.020 1.400 83.300 254.800 ;
      RECT 85.260 1.400 85.540 254.800 ;
      RECT 87.500 1.400 87.780 254.800 ;
      RECT 89.740 1.400 90.020 254.800 ;
      RECT 91.980 1.400 92.260 254.800 ;
      RECT 94.220 1.400 94.500 254.800 ;
      RECT 96.460 1.400 96.740 254.800 ;
      RECT 98.700 1.400 98.980 254.800 ;
      RECT 100.940 1.400 101.220 254.800 ;
      RECT 103.180 1.400 103.460 254.800 ;
      RECT 105.420 1.400 105.700 254.800 ;
      RECT 107.660 1.400 107.940 254.800 ;
      RECT 109.900 1.400 110.180 254.800 ;
      RECT 112.140 1.400 112.420 254.800 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 114.000 256.200 ;
    LAYER metal2 ;
    RECT 0 0 114.000 256.200 ;
    LAYER metal3 ;
    RECT 0.070 0 114.000 256.200 ;
    LAYER metal4 ;
    RECT 0 0 114.000 256.200 ;
    LAYER OVERLAP ;
    RECT 0 0 114.000 256.200 ;
  END
END liteeth_1rw1r_32w384d_8_sram

END LIBRARY
