VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_3x1_1r1w
  FOREIGN fakeram_3x1_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 70.110 BY 84.000 ;
  CLASS BLOCK ;
  PIN w_mask_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 -2.975 0.070 -2.905 ;
    END
  END w_mask_w1[0]
  PIN w_mask_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.505 0.070 1.575 ;
    END
  END w_mask_w1[1]
  PIN w_mask_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.985 0.070 6.055 ;
    END
  END w_mask_w1[2]
  PIN rd_out_r1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.125 0.070 6.195 ;
    END
  END rd_out_r1[0]
  PIN rd_out_r1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END rd_out_r1[1]
  PIN rd_out_r1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END rd_out_r1[2]
  PIN wd_in_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.225 0.070 15.295 ;
    END
  END wd_in_w1[0]
  PIN wd_in_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END wd_in_w1[1]
  PIN wd_in_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.185 0.070 24.255 ;
    END
  END wd_in_w1[2]
  PIN addr_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END addr_w1[0]
  PIN addr_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.805 0.070 28.875 ;
    END
  END addr_w1[1]
  PIN addr_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.285 0.070 33.355 ;
    END
  END addr_w1[2]
  PIN addr_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END addr_w1[3]
  PIN addr_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.245 0.070 42.315 ;
    END
  END addr_w1[4]
  PIN addr_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.725 0.070 46.795 ;
    END
  END addr_w1[5]
  PIN addr_r1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.865 0.070 46.935 ;
    END
  END addr_r1[0]
  PIN addr_r1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.345 0.070 51.415 ;
    END
  END addr_r1[1]
  PIN addr_r1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END addr_r1[2]
  PIN addr_r1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.305 0.070 60.375 ;
    END
  END addr_r1[3]
  PIN addr_r1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.785 0.070 64.855 ;
    END
  END addr_r1[4]
  PIN addr_r1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END addr_r1[5]
  PIN we_in_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.405 0.070 69.475 ;
    END
  END we_in_w1
  PIN ce_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.205 0.070 65.275 ;
    END
  END ce_w1
  PIN ce_r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.345 0.070 65.415 ;
    END
  END ce_r1
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.485 0.070 65.555 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 82.600 ;
      RECT 3.500 1.400 3.780 82.600 ;
      RECT 5.740 1.400 6.020 82.600 ;
      RECT 7.980 1.400 8.260 82.600 ;
      RECT 10.220 1.400 10.500 82.600 ;
      RECT 12.460 1.400 12.740 82.600 ;
      RECT 14.700 1.400 14.980 82.600 ;
      RECT 16.940 1.400 17.220 82.600 ;
      RECT 19.180 1.400 19.460 82.600 ;
      RECT 21.420 1.400 21.700 82.600 ;
      RECT 23.660 1.400 23.940 82.600 ;
      RECT 25.900 1.400 26.180 82.600 ;
      RECT 28.140 1.400 28.420 82.600 ;
      RECT 30.380 1.400 30.660 82.600 ;
      RECT 32.620 1.400 32.900 82.600 ;
      RECT 34.860 1.400 35.140 82.600 ;
      RECT 37.100 1.400 37.380 82.600 ;
      RECT 39.340 1.400 39.620 82.600 ;
      RECT 41.580 1.400 41.860 82.600 ;
      RECT 43.820 1.400 44.100 82.600 ;
      RECT 46.060 1.400 46.340 82.600 ;
      RECT 48.300 1.400 48.580 82.600 ;
      RECT 50.540 1.400 50.820 82.600 ;
      RECT 52.780 1.400 53.060 82.600 ;
      RECT 55.020 1.400 55.300 82.600 ;
      RECT 57.260 1.400 57.540 82.600 ;
      RECT 59.500 1.400 59.780 82.600 ;
      RECT 61.740 1.400 62.020 82.600 ;
      RECT 63.980 1.400 64.260 82.600 ;
      RECT 66.220 1.400 66.500 82.600 ;
      RECT 68.460 1.400 68.740 82.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 82.600 ;
      RECT 4.620 1.400 4.900 82.600 ;
      RECT 6.860 1.400 7.140 82.600 ;
      RECT 9.100 1.400 9.380 82.600 ;
      RECT 11.340 1.400 11.620 82.600 ;
      RECT 13.580 1.400 13.860 82.600 ;
      RECT 15.820 1.400 16.100 82.600 ;
      RECT 18.060 1.400 18.340 82.600 ;
      RECT 20.300 1.400 20.580 82.600 ;
      RECT 22.540 1.400 22.820 82.600 ;
      RECT 24.780 1.400 25.060 82.600 ;
      RECT 27.020 1.400 27.300 82.600 ;
      RECT 29.260 1.400 29.540 82.600 ;
      RECT 31.500 1.400 31.780 82.600 ;
      RECT 33.740 1.400 34.020 82.600 ;
      RECT 35.980 1.400 36.260 82.600 ;
      RECT 38.220 1.400 38.500 82.600 ;
      RECT 40.460 1.400 40.740 82.600 ;
      RECT 42.700 1.400 42.980 82.600 ;
      RECT 44.940 1.400 45.220 82.600 ;
      RECT 47.180 1.400 47.460 82.600 ;
      RECT 49.420 1.400 49.700 82.600 ;
      RECT 51.660 1.400 51.940 82.600 ;
      RECT 53.900 1.400 54.180 82.600 ;
      RECT 56.140 1.400 56.420 82.600 ;
      RECT 58.380 1.400 58.660 82.600 ;
      RECT 60.620 1.400 60.900 82.600 ;
      RECT 62.860 1.400 63.140 82.600 ;
      RECT 65.100 1.400 65.380 82.600 ;
      RECT 67.340 1.400 67.620 82.600 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 70.110 84.000 ;
    LAYER metal2 ;
    RECT 0 0 70.110 84.000 ;
    LAYER metal3 ;
    RECT 0.070 0 70.110 84.000 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 5.845 ;
    RECT 0 5.915 0.070 10.325 ;
    RECT 0 10.395 0.070 10.465 ;
    RECT 0 10.535 0.070 14.945 ;
    RECT 0 15.015 0.070 19.425 ;
    RECT 0 19.495 0.070 19.565 ;
    RECT 0 19.635 0.070 24.045 ;
    RECT 0 24.115 0.070 28.525 ;
    RECT 0 28.595 0.070 28.665 ;
    RECT 0 28.735 0.070 33.145 ;
    RECT 0 33.215 0.070 37.625 ;
    RECT 0 37.695 0.070 42.105 ;
    RECT 0 42.175 0.070 46.585 ;
    RECT 0 46.655 0.070 51.065 ;
    RECT 0 51.135 0.070 51.205 ;
    RECT 0 51.275 0.070 55.685 ;
    RECT 0 55.755 0.070 60.165 ;
    RECT 0 60.235 0.070 84.000 ;
    LAYER metal4 ;
    RECT 0 0 70.110 1.400 ;
    RECT 0 82.600 70.110 84.000 ;
    RECT 0.000 1.400 1.260 82.600 ;
    RECT 1.540 1.400 2.380 82.600 ;
    RECT 2.660 1.400 3.500 82.600 ;
    RECT 3.780 1.400 4.620 82.600 ;
    RECT 4.900 1.400 5.740 82.600 ;
    RECT 6.020 1.400 6.860 82.600 ;
    RECT 7.140 1.400 7.980 82.600 ;
    RECT 8.260 1.400 9.100 82.600 ;
    RECT 9.380 1.400 10.220 82.600 ;
    RECT 10.500 1.400 11.340 82.600 ;
    RECT 11.620 1.400 12.460 82.600 ;
    RECT 12.740 1.400 13.580 82.600 ;
    RECT 13.860 1.400 14.700 82.600 ;
    RECT 14.980 1.400 15.820 82.600 ;
    RECT 16.100 1.400 16.940 82.600 ;
    RECT 17.220 1.400 18.060 82.600 ;
    RECT 18.340 1.400 19.180 82.600 ;
    RECT 19.460 1.400 20.300 82.600 ;
    RECT 20.580 1.400 21.420 82.600 ;
    RECT 21.700 1.400 22.540 82.600 ;
    RECT 22.820 1.400 23.660 82.600 ;
    RECT 23.940 1.400 24.780 82.600 ;
    RECT 25.060 1.400 25.900 82.600 ;
    RECT 26.180 1.400 27.020 82.600 ;
    RECT 27.300 1.400 28.140 82.600 ;
    RECT 28.420 1.400 29.260 82.600 ;
    RECT 29.540 1.400 30.380 82.600 ;
    RECT 30.660 1.400 31.500 82.600 ;
    RECT 31.780 1.400 32.620 82.600 ;
    RECT 32.900 1.400 33.740 82.600 ;
    RECT 34.020 1.400 34.860 82.600 ;
    RECT 35.140 1.400 35.980 82.600 ;
    RECT 36.260 1.400 37.100 82.600 ;
    RECT 37.380 1.400 38.220 82.600 ;
    RECT 38.500 1.400 39.340 82.600 ;
    RECT 39.620 1.400 40.460 82.600 ;
    RECT 40.740 1.400 41.580 82.600 ;
    RECT 41.860 1.400 42.700 82.600 ;
    RECT 42.980 1.400 43.820 82.600 ;
    RECT 44.100 1.400 44.940 82.600 ;
    RECT 45.220 1.400 46.060 82.600 ;
    RECT 46.340 1.400 47.180 82.600 ;
    RECT 47.460 1.400 48.300 82.600 ;
    RECT 48.580 1.400 49.420 82.600 ;
    RECT 49.700 1.400 50.540 82.600 ;
    RECT 50.820 1.400 51.660 82.600 ;
    RECT 51.940 1.400 52.780 82.600 ;
    RECT 53.060 1.400 53.900 82.600 ;
    RECT 54.180 1.400 55.020 82.600 ;
    RECT 55.300 1.400 56.140 82.600 ;
    RECT 56.420 1.400 57.260 82.600 ;
    RECT 57.540 1.400 58.380 82.600 ;
    RECT 58.660 1.400 59.500 82.600 ;
    RECT 59.780 1.400 60.620 82.600 ;
    RECT 60.900 1.400 61.740 82.600 ;
    RECT 62.020 1.400 62.860 82.600 ;
    RECT 63.140 1.400 63.980 82.600 ;
    RECT 64.260 1.400 65.100 82.600 ;
    RECT 65.380 1.400 66.220 82.600 ;
    RECT 66.500 1.400 67.340 82.600 ;
    RECT 67.620 1.400 68.460 82.600 ;
    RECT 68.740 1.400 70.110 82.600 ;
    LAYER OVERLAP ;
    RECT 0 0 70.110 84.000 ;
  END
END fakeram_3x1_1r1w

END LIBRARY
