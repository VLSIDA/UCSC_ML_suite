VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_32x128_2r1w
  FOREIGN sram_32x128_2r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 96.710 BY 250.600 ;
  CLASS BLOCK ;
  PIN w_mask_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.645 0.070 1.715 ;
    END
  END w_mask_w1[0]
  PIN w_mask_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.885 0.070 3.955 ;
    END
  END w_mask_w1[1]
  PIN w_mask_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.125 0.070 6.195 ;
    END
  END w_mask_w1[2]
  PIN w_mask_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_w1[3]
  PIN w_mask_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_w1[4]
  PIN w_mask_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.845 0.070 12.915 ;
    END
  END w_mask_w1[5]
  PIN w_mask_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_w1[6]
  PIN w_mask_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.325 0.070 17.395 ;
    END
  END w_mask_w1[7]
  PIN w_mask_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.565 0.070 19.635 ;
    END
  END w_mask_w1[8]
  PIN w_mask_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_w1[9]
  PIN w_mask_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.045 0.070 24.115 ;
    END
  END w_mask_w1[10]
  PIN w_mask_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.285 0.070 26.355 ;
    END
  END w_mask_w1[11]
  PIN w_mask_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END w_mask_w1[12]
  PIN w_mask_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_w1[13]
  PIN w_mask_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.005 0.070 33.075 ;
    END
  END w_mask_w1[14]
  PIN w_mask_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END w_mask_w1[15]
  PIN w_mask_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.485 0.070 37.555 ;
    END
  END w_mask_w1[16]
  PIN w_mask_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.725 0.070 39.795 ;
    END
  END w_mask_w1[17]
  PIN w_mask_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END w_mask_w1[18]
  PIN w_mask_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.205 0.070 44.275 ;
    END
  END w_mask_w1[19]
  PIN w_mask_w1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.445 0.070 46.515 ;
    END
  END w_mask_w1[20]
  PIN w_mask_w1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END w_mask_w1[21]
  PIN w_mask_w1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.925 0.070 50.995 ;
    END
  END w_mask_w1[22]
  PIN w_mask_w1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.165 0.070 53.235 ;
    END
  END w_mask_w1[23]
  PIN w_mask_w1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END w_mask_w1[24]
  PIN w_mask_w1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.645 0.070 57.715 ;
    END
  END w_mask_w1[25]
  PIN w_mask_w1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.885 0.070 59.955 ;
    END
  END w_mask_w1[26]
  PIN w_mask_w1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END w_mask_w1[27]
  PIN w_mask_w1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.365 0.070 64.435 ;
    END
  END w_mask_w1[28]
  PIN w_mask_w1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.605 0.070 66.675 ;
    END
  END w_mask_w1[29]
  PIN w_mask_w1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END w_mask_w1[30]
  PIN w_mask_w1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.085 0.070 71.155 ;
    END
  END w_mask_w1[31]
  PIN rd_out_r1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.605 0.070 73.675 ;
    END
  END rd_out_r1[0]
  PIN rd_out_r1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.845 0.070 75.915 ;
    END
  END rd_out_r1[1]
  PIN rd_out_r1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END rd_out_r1[2]
  PIN rd_out_r1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.325 0.070 80.395 ;
    END
  END rd_out_r1[3]
  PIN rd_out_r1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.565 0.070 82.635 ;
    END
  END rd_out_r1[4]
  PIN rd_out_r1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END rd_out_r1[5]
  PIN rd_out_r1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.045 0.070 87.115 ;
    END
  END rd_out_r1[6]
  PIN rd_out_r1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.285 0.070 89.355 ;
    END
  END rd_out_r1[7]
  PIN rd_out_r1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END rd_out_r1[8]
  PIN rd_out_r1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.765 0.070 93.835 ;
    END
  END rd_out_r1[9]
  PIN rd_out_r1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.005 0.070 96.075 ;
    END
  END rd_out_r1[10]
  PIN rd_out_r1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.245 0.070 98.315 ;
    END
  END rd_out_r1[11]
  PIN rd_out_r1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.485 0.070 100.555 ;
    END
  END rd_out_r1[12]
  PIN rd_out_r1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.725 0.070 102.795 ;
    END
  END rd_out_r1[13]
  PIN rd_out_r1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.965 0.070 105.035 ;
    END
  END rd_out_r1[14]
  PIN rd_out_r1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.205 0.070 107.275 ;
    END
  END rd_out_r1[15]
  PIN rd_out_r1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.445 0.070 109.515 ;
    END
  END rd_out_r1[16]
  PIN rd_out_r1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.685 0.070 111.755 ;
    END
  END rd_out_r1[17]
  PIN rd_out_r1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.925 0.070 113.995 ;
    END
  END rd_out_r1[18]
  PIN rd_out_r1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.165 0.070 116.235 ;
    END
  END rd_out_r1[19]
  PIN rd_out_r1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.405 0.070 118.475 ;
    END
  END rd_out_r1[20]
  PIN rd_out_r1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.645 0.070 120.715 ;
    END
  END rd_out_r1[21]
  PIN rd_out_r1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.885 0.070 122.955 ;
    END
  END rd_out_r1[22]
  PIN rd_out_r1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.125 0.070 125.195 ;
    END
  END rd_out_r1[23]
  PIN rd_out_r1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.365 0.070 127.435 ;
    END
  END rd_out_r1[24]
  PIN rd_out_r1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.605 0.070 129.675 ;
    END
  END rd_out_r1[25]
  PIN rd_out_r1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.845 0.070 131.915 ;
    END
  END rd_out_r1[26]
  PIN rd_out_r1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.085 0.070 134.155 ;
    END
  END rd_out_r1[27]
  PIN rd_out_r1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.325 0.070 136.395 ;
    END
  END rd_out_r1[28]
  PIN rd_out_r1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.565 0.070 138.635 ;
    END
  END rd_out_r1[29]
  PIN rd_out_r1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.805 0.070 140.875 ;
    END
  END rd_out_r1[30]
  PIN rd_out_r1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.045 0.070 143.115 ;
    END
  END rd_out_r1[31]
  PIN rd_out_r2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.565 0.070 145.635 ;
    END
  END rd_out_r2[0]
  PIN rd_out_r2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.805 0.070 147.875 ;
    END
  END rd_out_r2[1]
  PIN rd_out_r2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.045 0.070 150.115 ;
    END
  END rd_out_r2[2]
  PIN rd_out_r2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.285 0.070 152.355 ;
    END
  END rd_out_r2[3]
  PIN rd_out_r2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.525 0.070 154.595 ;
    END
  END rd_out_r2[4]
  PIN rd_out_r2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.765 0.070 156.835 ;
    END
  END rd_out_r2[5]
  PIN rd_out_r2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.005 0.070 159.075 ;
    END
  END rd_out_r2[6]
  PIN rd_out_r2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.245 0.070 161.315 ;
    END
  END rd_out_r2[7]
  PIN rd_out_r2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.485 0.070 163.555 ;
    END
  END rd_out_r2[8]
  PIN rd_out_r2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.725 0.070 165.795 ;
    END
  END rd_out_r2[9]
  PIN rd_out_r2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.965 0.070 168.035 ;
    END
  END rd_out_r2[10]
  PIN rd_out_r2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.205 0.070 170.275 ;
    END
  END rd_out_r2[11]
  PIN rd_out_r2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.445 0.070 172.515 ;
    END
  END rd_out_r2[12]
  PIN rd_out_r2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.685 0.070 174.755 ;
    END
  END rd_out_r2[13]
  PIN rd_out_r2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.925 0.070 176.995 ;
    END
  END rd_out_r2[14]
  PIN rd_out_r2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.165 0.070 179.235 ;
    END
  END rd_out_r2[15]
  PIN rd_out_r2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.405 0.070 181.475 ;
    END
  END rd_out_r2[16]
  PIN rd_out_r2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.645 0.070 183.715 ;
    END
  END rd_out_r2[17]
  PIN rd_out_r2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.885 0.070 185.955 ;
    END
  END rd_out_r2[18]
  PIN rd_out_r2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.125 0.070 188.195 ;
    END
  END rd_out_r2[19]
  PIN rd_out_r2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.365 0.070 190.435 ;
    END
  END rd_out_r2[20]
  PIN rd_out_r2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.605 0.070 192.675 ;
    END
  END rd_out_r2[21]
  PIN rd_out_r2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.845 0.070 194.915 ;
    END
  END rd_out_r2[22]
  PIN rd_out_r2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.085 0.070 197.155 ;
    END
  END rd_out_r2[23]
  PIN rd_out_r2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.325 0.070 199.395 ;
    END
  END rd_out_r2[24]
  PIN rd_out_r2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.565 0.070 201.635 ;
    END
  END rd_out_r2[25]
  PIN rd_out_r2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.805 0.070 203.875 ;
    END
  END rd_out_r2[26]
  PIN rd_out_r2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.045 0.070 206.115 ;
    END
  END rd_out_r2[27]
  PIN rd_out_r2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.285 0.070 208.355 ;
    END
  END rd_out_r2[28]
  PIN rd_out_r2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.525 0.070 210.595 ;
    END
  END rd_out_r2[29]
  PIN rd_out_r2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.765 0.070 212.835 ;
    END
  END rd_out_r2[30]
  PIN rd_out_r2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.005 0.070 215.075 ;
    END
  END rd_out_r2[31]
  PIN wd_in_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.525 0.070 217.595 ;
    END
  END wd_in_w1[0]
  PIN wd_in_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.765 0.070 219.835 ;
    END
  END wd_in_w1[1]
  PIN wd_in_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.005 0.070 222.075 ;
    END
  END wd_in_w1[2]
  PIN wd_in_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.245 0.070 224.315 ;
    END
  END wd_in_w1[3]
  PIN wd_in_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.485 0.070 226.555 ;
    END
  END wd_in_w1[4]
  PIN wd_in_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.725 0.070 228.795 ;
    END
  END wd_in_w1[5]
  PIN wd_in_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.965 0.070 231.035 ;
    END
  END wd_in_w1[6]
  PIN wd_in_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.205 0.070 233.275 ;
    END
  END wd_in_w1[7]
  PIN wd_in_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.445 0.070 235.515 ;
    END
  END wd_in_w1[8]
  PIN wd_in_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.685 0.070 237.755 ;
    END
  END wd_in_w1[9]
  PIN wd_in_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.925 0.070 239.995 ;
    END
  END wd_in_w1[10]
  PIN wd_in_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.165 0.070 242.235 ;
    END
  END wd_in_w1[11]
  PIN wd_in_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.405 0.070 244.475 ;
    END
  END wd_in_w1[12]
  PIN wd_in_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.645 0.070 246.715 ;
    END
  END wd_in_w1[13]
  PIN wd_in_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.885 0.070 248.955 ;
    END
  END wd_in_w1[14]
  PIN wd_in_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.125 0.070 251.195 ;
    END
  END wd_in_w1[15]
  PIN wd_in_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.365 0.070 253.435 ;
    END
  END wd_in_w1[16]
  PIN wd_in_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.605 0.070 255.675 ;
    END
  END wd_in_w1[17]
  PIN wd_in_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.845 0.070 257.915 ;
    END
  END wd_in_w1[18]
  PIN wd_in_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.085 0.070 260.155 ;
    END
  END wd_in_w1[19]
  PIN wd_in_w1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.325 0.070 262.395 ;
    END
  END wd_in_w1[20]
  PIN wd_in_w1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.565 0.070 264.635 ;
    END
  END wd_in_w1[21]
  PIN wd_in_w1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.805 0.070 266.875 ;
    END
  END wd_in_w1[22]
  PIN wd_in_w1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.045 0.070 269.115 ;
    END
  END wd_in_w1[23]
  PIN wd_in_w1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.285 0.070 271.355 ;
    END
  END wd_in_w1[24]
  PIN wd_in_w1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.525 0.070 273.595 ;
    END
  END wd_in_w1[25]
  PIN wd_in_w1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.765 0.070 275.835 ;
    END
  END wd_in_w1[26]
  PIN wd_in_w1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.005 0.070 278.075 ;
    END
  END wd_in_w1[27]
  PIN wd_in_w1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.245 0.070 280.315 ;
    END
  END wd_in_w1[28]
  PIN wd_in_w1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.485 0.070 282.555 ;
    END
  END wd_in_w1[29]
  PIN wd_in_w1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.725 0.070 284.795 ;
    END
  END wd_in_w1[30]
  PIN wd_in_w1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.965 0.070 287.035 ;
    END
  END wd_in_w1[31]
  PIN addr_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.485 0.070 289.555 ;
    END
  END addr_w1[0]
  PIN addr_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.725 0.070 291.795 ;
    END
  END addr_w1[1]
  PIN addr_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.965 0.070 294.035 ;
    END
  END addr_w1[2]
  PIN addr_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.205 0.070 296.275 ;
    END
  END addr_w1[3]
  PIN addr_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.445 0.070 298.515 ;
    END
  END addr_w1[4]
  PIN addr_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.685 0.070 300.755 ;
    END
  END addr_w1[5]
  PIN addr_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.925 0.070 302.995 ;
    END
  END addr_w1[6]
  PIN addr_r1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.445 0.070 305.515 ;
    END
  END addr_r1[0]
  PIN addr_r1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.685 0.070 307.755 ;
    END
  END addr_r1[1]
  PIN addr_r1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.925 0.070 309.995 ;
    END
  END addr_r1[2]
  PIN addr_r1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.165 0.070 312.235 ;
    END
  END addr_r1[3]
  PIN addr_r1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.405 0.070 314.475 ;
    END
  END addr_r1[4]
  PIN addr_r1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.645 0.070 316.715 ;
    END
  END addr_r1[5]
  PIN addr_r1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.885 0.070 318.955 ;
    END
  END addr_r1[6]
  PIN addr_r2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.405 0.070 321.475 ;
    END
  END addr_r2[0]
  PIN addr_r2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.645 0.070 323.715 ;
    END
  END addr_r2[1]
  PIN addr_r2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.885 0.070 325.955 ;
    END
  END addr_r2[2]
  PIN addr_r2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.125 0.070 328.195 ;
    END
  END addr_r2[3]
  PIN addr_r2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 330.365 0.070 330.435 ;
    END
  END addr_r2[4]
  PIN addr_r2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.605 0.070 332.675 ;
    END
  END addr_r2[5]
  PIN addr_r2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.845 0.070 334.915 ;
    END
  END addr_r2[6]
  PIN we_in_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.365 0.070 337.435 ;
    END
  END we_in_w1
  PIN ce_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.165 0.070 340.235 ;
    END
  END ce_w1
  PIN ce_r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.685 0.070 342.755 ;
    END
  END ce_r1
  PIN ce_r2
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.925 0.070 344.995 ;
    END
  END ce_r2
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.445 0.070 347.515 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 249.200 ;
      RECT 3.500 1.400 3.780 249.200 ;
      RECT 5.740 1.400 6.020 249.200 ;
      RECT 7.980 1.400 8.260 249.200 ;
      RECT 10.220 1.400 10.500 249.200 ;
      RECT 12.460 1.400 12.740 249.200 ;
      RECT 14.700 1.400 14.980 249.200 ;
      RECT 16.940 1.400 17.220 249.200 ;
      RECT 19.180 1.400 19.460 249.200 ;
      RECT 21.420 1.400 21.700 249.200 ;
      RECT 23.660 1.400 23.940 249.200 ;
      RECT 25.900 1.400 26.180 249.200 ;
      RECT 28.140 1.400 28.420 249.200 ;
      RECT 30.380 1.400 30.660 249.200 ;
      RECT 32.620 1.400 32.900 249.200 ;
      RECT 34.860 1.400 35.140 249.200 ;
      RECT 37.100 1.400 37.380 249.200 ;
      RECT 39.340 1.400 39.620 249.200 ;
      RECT 41.580 1.400 41.860 249.200 ;
      RECT 43.820 1.400 44.100 249.200 ;
      RECT 46.060 1.400 46.340 249.200 ;
      RECT 48.300 1.400 48.580 249.200 ;
      RECT 50.540 1.400 50.820 249.200 ;
      RECT 52.780 1.400 53.060 249.200 ;
      RECT 55.020 1.400 55.300 249.200 ;
      RECT 57.260 1.400 57.540 249.200 ;
      RECT 59.500 1.400 59.780 249.200 ;
      RECT 61.740 1.400 62.020 249.200 ;
      RECT 63.980 1.400 64.260 249.200 ;
      RECT 66.220 1.400 66.500 249.200 ;
      RECT 68.460 1.400 68.740 249.200 ;
      RECT 70.700 1.400 70.980 249.200 ;
      RECT 72.940 1.400 73.220 249.200 ;
      RECT 75.180 1.400 75.460 249.200 ;
      RECT 77.420 1.400 77.700 249.200 ;
      RECT 79.660 1.400 79.940 249.200 ;
      RECT 81.900 1.400 82.180 249.200 ;
      RECT 84.140 1.400 84.420 249.200 ;
      RECT 86.380 1.400 86.660 249.200 ;
      RECT 88.620 1.400 88.900 249.200 ;
      RECT 90.860 1.400 91.140 249.200 ;
      RECT 93.100 1.400 93.380 249.200 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 249.200 ;
      RECT 4.620 1.400 4.900 249.200 ;
      RECT 6.860 1.400 7.140 249.200 ;
      RECT 9.100 1.400 9.380 249.200 ;
      RECT 11.340 1.400 11.620 249.200 ;
      RECT 13.580 1.400 13.860 249.200 ;
      RECT 15.820 1.400 16.100 249.200 ;
      RECT 18.060 1.400 18.340 249.200 ;
      RECT 20.300 1.400 20.580 249.200 ;
      RECT 22.540 1.400 22.820 249.200 ;
      RECT 24.780 1.400 25.060 249.200 ;
      RECT 27.020 1.400 27.300 249.200 ;
      RECT 29.260 1.400 29.540 249.200 ;
      RECT 31.500 1.400 31.780 249.200 ;
      RECT 33.740 1.400 34.020 249.200 ;
      RECT 35.980 1.400 36.260 249.200 ;
      RECT 38.220 1.400 38.500 249.200 ;
      RECT 40.460 1.400 40.740 249.200 ;
      RECT 42.700 1.400 42.980 249.200 ;
      RECT 44.940 1.400 45.220 249.200 ;
      RECT 47.180 1.400 47.460 249.200 ;
      RECT 49.420 1.400 49.700 249.200 ;
      RECT 51.660 1.400 51.940 249.200 ;
      RECT 53.900 1.400 54.180 249.200 ;
      RECT 56.140 1.400 56.420 249.200 ;
      RECT 58.380 1.400 58.660 249.200 ;
      RECT 60.620 1.400 60.900 249.200 ;
      RECT 62.860 1.400 63.140 249.200 ;
      RECT 65.100 1.400 65.380 249.200 ;
      RECT 67.340 1.400 67.620 249.200 ;
      RECT 69.580 1.400 69.860 249.200 ;
      RECT 71.820 1.400 72.100 249.200 ;
      RECT 74.060 1.400 74.340 249.200 ;
      RECT 76.300 1.400 76.580 249.200 ;
      RECT 78.540 1.400 78.820 249.200 ;
      RECT 80.780 1.400 81.060 249.200 ;
      RECT 83.020 1.400 83.300 249.200 ;
      RECT 85.260 1.400 85.540 249.200 ;
      RECT 87.500 1.400 87.780 249.200 ;
      RECT 89.740 1.400 90.020 249.200 ;
      RECT 91.980 1.400 92.260 249.200 ;
      RECT 94.220 1.400 94.500 249.200 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 96.710 250.600 ;
    LAYER metal2 ;
    RECT 0 0 96.710 250.600 ;
    LAYER metal3 ;
    RECT 0.070 0 96.710 250.600 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 3.605 ;
    RECT 0 3.675 0.070 5.845 ;
    RECT 0 5.915 0.070 8.085 ;
    RECT 0 8.155 0.070 10.325 ;
    RECT 0 10.395 0.070 12.565 ;
    RECT 0 12.635 0.070 14.805 ;
    RECT 0 14.875 0.070 17.045 ;
    RECT 0 17.115 0.070 19.285 ;
    RECT 0 19.355 0.070 21.525 ;
    RECT 0 21.595 0.070 23.765 ;
    RECT 0 23.835 0.070 26.005 ;
    RECT 0 26.075 0.070 28.245 ;
    RECT 0 28.315 0.070 30.485 ;
    RECT 0 30.555 0.070 32.725 ;
    RECT 0 32.795 0.070 34.965 ;
    RECT 0 35.035 0.070 37.205 ;
    RECT 0 37.275 0.070 39.445 ;
    RECT 0 39.515 0.070 41.685 ;
    RECT 0 41.755 0.070 43.925 ;
    RECT 0 43.995 0.070 46.165 ;
    RECT 0 46.235 0.070 48.405 ;
    RECT 0 48.475 0.070 50.645 ;
    RECT 0 50.715 0.070 52.885 ;
    RECT 0 52.955 0.070 55.125 ;
    RECT 0 55.195 0.070 57.365 ;
    RECT 0 57.435 0.070 59.605 ;
    RECT 0 59.675 0.070 61.845 ;
    RECT 0 61.915 0.070 64.085 ;
    RECT 0 64.155 0.070 66.325 ;
    RECT 0 66.395 0.070 68.565 ;
    RECT 0 68.635 0.070 70.805 ;
    RECT 0 70.875 0.070 73.325 ;
    RECT 0 73.395 0.070 75.565 ;
    RECT 0 75.635 0.070 77.805 ;
    RECT 0 77.875 0.070 80.045 ;
    RECT 0 80.115 0.070 82.285 ;
    RECT 0 82.355 0.070 84.525 ;
    RECT 0 84.595 0.070 86.765 ;
    RECT 0 86.835 0.070 89.005 ;
    RECT 0 89.075 0.070 91.245 ;
    RECT 0 91.315 0.070 93.485 ;
    RECT 0 93.555 0.070 95.725 ;
    RECT 0 95.795 0.070 97.965 ;
    RECT 0 98.035 0.070 100.205 ;
    RECT 0 100.275 0.070 102.445 ;
    RECT 0 102.515 0.070 104.685 ;
    RECT 0 104.755 0.070 106.925 ;
    RECT 0 106.995 0.070 109.165 ;
    RECT 0 109.235 0.070 111.405 ;
    RECT 0 111.475 0.070 113.645 ;
    RECT 0 113.715 0.070 115.885 ;
    RECT 0 115.955 0.070 118.125 ;
    RECT 0 118.195 0.070 120.365 ;
    RECT 0 120.435 0.070 122.605 ;
    RECT 0 122.675 0.070 124.845 ;
    RECT 0 124.915 0.070 127.085 ;
    RECT 0 127.155 0.070 129.325 ;
    RECT 0 129.395 0.070 131.565 ;
    RECT 0 131.635 0.070 133.805 ;
    RECT 0 133.875 0.070 136.045 ;
    RECT 0 136.115 0.070 138.285 ;
    RECT 0 138.355 0.070 140.525 ;
    RECT 0 140.595 0.070 142.765 ;
    RECT 0 142.835 0.070 145.285 ;
    RECT 0 145.355 0.070 147.525 ;
    RECT 0 147.595 0.070 149.765 ;
    RECT 0 149.835 0.070 152.005 ;
    RECT 0 152.075 0.070 154.245 ;
    RECT 0 154.315 0.070 156.485 ;
    RECT 0 156.555 0.070 158.725 ;
    RECT 0 158.795 0.070 160.965 ;
    RECT 0 161.035 0.070 163.205 ;
    RECT 0 163.275 0.070 165.445 ;
    RECT 0 165.515 0.070 167.685 ;
    RECT 0 167.755 0.070 169.925 ;
    RECT 0 169.995 0.070 172.165 ;
    RECT 0 172.235 0.070 174.405 ;
    RECT 0 174.475 0.070 176.645 ;
    RECT 0 176.715 0.070 178.885 ;
    RECT 0 178.955 0.070 181.125 ;
    RECT 0 181.195 0.070 183.365 ;
    RECT 0 183.435 0.070 185.605 ;
    RECT 0 185.675 0.070 187.845 ;
    RECT 0 187.915 0.070 190.085 ;
    RECT 0 190.155 0.070 192.325 ;
    RECT 0 192.395 0.070 194.565 ;
    RECT 0 194.635 0.070 196.805 ;
    RECT 0 196.875 0.070 199.045 ;
    RECT 0 199.115 0.070 201.285 ;
    RECT 0 201.355 0.070 203.525 ;
    RECT 0 203.595 0.070 205.765 ;
    RECT 0 205.835 0.070 208.005 ;
    RECT 0 208.075 0.070 210.245 ;
    RECT 0 210.315 0.070 212.485 ;
    RECT 0 212.555 0.070 214.725 ;
    RECT 0 214.795 0.070 217.245 ;
    RECT 0 217.315 0.070 219.485 ;
    RECT 0 219.555 0.070 221.725 ;
    RECT 0 221.795 0.070 223.965 ;
    RECT 0 224.035 0.070 226.205 ;
    RECT 0 226.275 0.070 228.445 ;
    RECT 0 228.515 0.070 230.685 ;
    RECT 0 230.755 0.070 233.205 ;
    RECT 0 233.275 0.070 235.445 ;
    RECT 0 235.515 0.070 237.685 ;
    RECT 0 237.755 0.070 250.600 ;
    LAYER metal4 ;
    RECT 0 0 96.710 1.400 ;
    RECT 0 249.200 96.710 250.600 ;
    RECT 0.000 1.400 1.260 249.200 ;
    RECT 1.540 1.400 2.380 249.200 ;
    RECT 2.660 1.400 3.500 249.200 ;
    RECT 3.780 1.400 4.620 249.200 ;
    RECT 4.900 1.400 5.740 249.200 ;
    RECT 6.020 1.400 6.860 249.200 ;
    RECT 7.140 1.400 7.980 249.200 ;
    RECT 8.260 1.400 9.100 249.200 ;
    RECT 9.380 1.400 10.220 249.200 ;
    RECT 10.500 1.400 11.340 249.200 ;
    RECT 11.620 1.400 12.460 249.200 ;
    RECT 12.740 1.400 13.580 249.200 ;
    RECT 13.860 1.400 14.700 249.200 ;
    RECT 14.980 1.400 15.820 249.200 ;
    RECT 16.100 1.400 16.940 249.200 ;
    RECT 17.220 1.400 18.060 249.200 ;
    RECT 18.340 1.400 19.180 249.200 ;
    RECT 19.460 1.400 20.300 249.200 ;
    RECT 20.580 1.400 21.420 249.200 ;
    RECT 21.700 1.400 22.540 249.200 ;
    RECT 22.820 1.400 23.660 249.200 ;
    RECT 23.940 1.400 24.780 249.200 ;
    RECT 25.060 1.400 25.900 249.200 ;
    RECT 26.180 1.400 27.020 249.200 ;
    RECT 27.300 1.400 28.140 249.200 ;
    RECT 28.420 1.400 29.260 249.200 ;
    RECT 29.540 1.400 30.380 249.200 ;
    RECT 30.660 1.400 31.500 249.200 ;
    RECT 31.780 1.400 32.620 249.200 ;
    RECT 32.900 1.400 33.740 249.200 ;
    RECT 34.020 1.400 34.860 249.200 ;
    RECT 35.140 1.400 35.980 249.200 ;
    RECT 36.260 1.400 37.100 249.200 ;
    RECT 37.380 1.400 38.220 249.200 ;
    RECT 38.500 1.400 39.340 249.200 ;
    RECT 39.620 1.400 40.460 249.200 ;
    RECT 40.740 1.400 41.580 249.200 ;
    RECT 41.860 1.400 42.700 249.200 ;
    RECT 42.980 1.400 43.820 249.200 ;
    RECT 44.100 1.400 44.940 249.200 ;
    RECT 45.220 1.400 46.060 249.200 ;
    RECT 46.340 1.400 47.180 249.200 ;
    RECT 47.460 1.400 48.300 249.200 ;
    RECT 48.580 1.400 49.420 249.200 ;
    RECT 49.700 1.400 50.540 249.200 ;
    RECT 50.820 1.400 51.660 249.200 ;
    RECT 51.940 1.400 52.780 249.200 ;
    RECT 53.060 1.400 53.900 249.200 ;
    RECT 54.180 1.400 55.020 249.200 ;
    RECT 55.300 1.400 56.140 249.200 ;
    RECT 56.420 1.400 57.260 249.200 ;
    RECT 57.540 1.400 58.380 249.200 ;
    RECT 58.660 1.400 59.500 249.200 ;
    RECT 59.780 1.400 60.620 249.200 ;
    RECT 60.900 1.400 61.740 249.200 ;
    RECT 62.020 1.400 62.860 249.200 ;
    RECT 63.140 1.400 63.980 249.200 ;
    RECT 64.260 1.400 65.100 249.200 ;
    RECT 65.380 1.400 66.220 249.200 ;
    RECT 66.500 1.400 67.340 249.200 ;
    RECT 67.620 1.400 68.460 249.200 ;
    RECT 68.740 1.400 69.580 249.200 ;
    RECT 69.860 1.400 70.700 249.200 ;
    RECT 70.980 1.400 71.820 249.200 ;
    RECT 72.100 1.400 72.940 249.200 ;
    RECT 73.220 1.400 74.060 249.200 ;
    RECT 74.340 1.400 75.180 249.200 ;
    RECT 75.460 1.400 76.300 249.200 ;
    RECT 76.580 1.400 77.420 249.200 ;
    RECT 77.700 1.400 78.540 249.200 ;
    RECT 78.820 1.400 79.660 249.200 ;
    RECT 79.940 1.400 80.780 249.200 ;
    RECT 81.060 1.400 81.900 249.200 ;
    RECT 82.180 1.400 83.020 249.200 ;
    RECT 83.300 1.400 84.140 249.200 ;
    RECT 84.420 1.400 85.260 249.200 ;
    RECT 85.540 1.400 86.380 249.200 ;
    RECT 86.660 1.400 87.500 249.200 ;
    RECT 87.780 1.400 88.620 249.200 ;
    RECT 88.900 1.400 89.740 249.200 ;
    RECT 90.020 1.400 90.860 249.200 ;
    RECT 91.140 1.400 91.980 249.200 ;
    RECT 92.260 1.400 93.100 249.200 ;
    RECT 93.380 1.400 94.220 249.200 ;
    RECT 94.500 1.400 96.710 249.200 ;
    LAYER OVERLAP ;
    RECT 0 0 96.710 250.600 ;
  END
END sram_32x128_2r1w

END LIBRARY
