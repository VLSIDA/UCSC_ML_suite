VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_512x256_1r1w
  FOREIGN fakeram_512x256_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 689.130 BY 767.200 ;
  CLASS BLOCK ;
  PIN w_mask_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.505 0.070 29.575 ;
    END
  END w_mask_w1[0]
  PIN w_mask_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.925 0.070 29.995 ;
    END
  END w_mask_w1[1]
  PIN w_mask_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.345 0.070 30.415 ;
    END
  END w_mask_w1[2]
  PIN w_mask_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_w1[3]
  PIN w_mask_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.185 0.070 31.255 ;
    END
  END w_mask_w1[4]
  PIN w_mask_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.605 0.070 31.675 ;
    END
  END w_mask_w1[5]
  PIN w_mask_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.025 0.070 32.095 ;
    END
  END w_mask_w1[6]
  PIN w_mask_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.445 0.070 32.515 ;
    END
  END w_mask_w1[7]
  PIN w_mask_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.865 0.070 32.935 ;
    END
  END w_mask_w1[8]
  PIN w_mask_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.285 0.070 33.355 ;
    END
  END w_mask_w1[9]
  PIN w_mask_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.705 0.070 33.775 ;
    END
  END w_mask_w1[10]
  PIN w_mask_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.125 0.070 34.195 ;
    END
  END w_mask_w1[11]
  PIN w_mask_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.545 0.070 34.615 ;
    END
  END w_mask_w1[12]
  PIN w_mask_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_w1[13]
  PIN w_mask_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.385 0.070 35.455 ;
    END
  END w_mask_w1[14]
  PIN w_mask_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.805 0.070 35.875 ;
    END
  END w_mask_w1[15]
  PIN w_mask_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.225 0.070 36.295 ;
    END
  END w_mask_w1[16]
  PIN w_mask_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END w_mask_w1[17]
  PIN w_mask_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.065 0.070 37.135 ;
    END
  END w_mask_w1[18]
  PIN w_mask_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.485 0.070 37.555 ;
    END
  END w_mask_w1[19]
  PIN w_mask_w1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.905 0.070 37.975 ;
    END
  END w_mask_w1[20]
  PIN w_mask_w1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.325 0.070 38.395 ;
    END
  END w_mask_w1[21]
  PIN w_mask_w1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.745 0.070 38.815 ;
    END
  END w_mask_w1[22]
  PIN w_mask_w1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END w_mask_w1[23]
  PIN w_mask_w1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.585 0.070 39.655 ;
    END
  END w_mask_w1[24]
  PIN w_mask_w1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.005 0.070 40.075 ;
    END
  END w_mask_w1[25]
  PIN w_mask_w1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.425 0.070 40.495 ;
    END
  END w_mask_w1[26]
  PIN w_mask_w1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.845 0.070 40.915 ;
    END
  END w_mask_w1[27]
  PIN w_mask_w1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.265 0.070 41.335 ;
    END
  END w_mask_w1[28]
  PIN w_mask_w1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.685 0.070 41.755 ;
    END
  END w_mask_w1[29]
  PIN w_mask_w1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.105 0.070 42.175 ;
    END
  END w_mask_w1[30]
  PIN w_mask_w1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END w_mask_w1[31]
  PIN w_mask_w1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.945 0.070 43.015 ;
    END
  END w_mask_w1[32]
  PIN w_mask_w1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END w_mask_w1[33]
  PIN w_mask_w1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.785 0.070 43.855 ;
    END
  END w_mask_w1[34]
  PIN w_mask_w1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.205 0.070 44.275 ;
    END
  END w_mask_w1[35]
  PIN w_mask_w1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.625 0.070 44.695 ;
    END
  END w_mask_w1[36]
  PIN w_mask_w1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END w_mask_w1[37]
  PIN w_mask_w1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.465 0.070 45.535 ;
    END
  END w_mask_w1[38]
  PIN w_mask_w1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.885 0.070 45.955 ;
    END
  END w_mask_w1[39]
  PIN w_mask_w1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.305 0.070 46.375 ;
    END
  END w_mask_w1[40]
  PIN w_mask_w1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.725 0.070 46.795 ;
    END
  END w_mask_w1[41]
  PIN w_mask_w1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.145 0.070 47.215 ;
    END
  END w_mask_w1[42]
  PIN w_mask_w1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.565 0.070 47.635 ;
    END
  END w_mask_w1[43]
  PIN w_mask_w1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.985 0.070 48.055 ;
    END
  END w_mask_w1[44]
  PIN w_mask_w1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END w_mask_w1[45]
  PIN w_mask_w1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.825 0.070 48.895 ;
    END
  END w_mask_w1[46]
  PIN w_mask_w1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.245 0.070 49.315 ;
    END
  END w_mask_w1[47]
  PIN w_mask_w1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.665 0.070 49.735 ;
    END
  END w_mask_w1[48]
  PIN w_mask_w1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.085 0.070 50.155 ;
    END
  END w_mask_w1[49]
  PIN w_mask_w1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.505 0.070 50.575 ;
    END
  END w_mask_w1[50]
  PIN w_mask_w1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.925 0.070 50.995 ;
    END
  END w_mask_w1[51]
  PIN w_mask_w1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.345 0.070 51.415 ;
    END
  END w_mask_w1[52]
  PIN w_mask_w1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.765 0.070 51.835 ;
    END
  END w_mask_w1[53]
  PIN w_mask_w1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.185 0.070 52.255 ;
    END
  END w_mask_w1[54]
  PIN w_mask_w1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.605 0.070 52.675 ;
    END
  END w_mask_w1[55]
  PIN w_mask_w1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.025 0.070 53.095 ;
    END
  END w_mask_w1[56]
  PIN w_mask_w1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.445 0.070 53.515 ;
    END
  END w_mask_w1[57]
  PIN w_mask_w1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.865 0.070 53.935 ;
    END
  END w_mask_w1[58]
  PIN w_mask_w1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.285 0.070 54.355 ;
    END
  END w_mask_w1[59]
  PIN w_mask_w1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.705 0.070 54.775 ;
    END
  END w_mask_w1[60]
  PIN w_mask_w1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.125 0.070 55.195 ;
    END
  END w_mask_w1[61]
  PIN w_mask_w1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.545 0.070 55.615 ;
    END
  END w_mask_w1[62]
  PIN w_mask_w1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.965 0.070 56.035 ;
    END
  END w_mask_w1[63]
  PIN w_mask_w1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.385 0.070 56.455 ;
    END
  END w_mask_w1[64]
  PIN w_mask_w1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.805 0.070 56.875 ;
    END
  END w_mask_w1[65]
  PIN w_mask_w1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.225 0.070 57.295 ;
    END
  END w_mask_w1[66]
  PIN w_mask_w1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.645 0.070 57.715 ;
    END
  END w_mask_w1[67]
  PIN w_mask_w1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.065 0.070 58.135 ;
    END
  END w_mask_w1[68]
  PIN w_mask_w1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.485 0.070 58.555 ;
    END
  END w_mask_w1[69]
  PIN w_mask_w1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.905 0.070 58.975 ;
    END
  END w_mask_w1[70]
  PIN w_mask_w1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.325 0.070 59.395 ;
    END
  END w_mask_w1[71]
  PIN w_mask_w1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.745 0.070 59.815 ;
    END
  END w_mask_w1[72]
  PIN w_mask_w1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_w1[73]
  PIN w_mask_w1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.585 0.070 60.655 ;
    END
  END w_mask_w1[74]
  PIN w_mask_w1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.005 0.070 61.075 ;
    END
  END w_mask_w1[75]
  PIN w_mask_w1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.425 0.070 61.495 ;
    END
  END w_mask_w1[76]
  PIN w_mask_w1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.845 0.070 61.915 ;
    END
  END w_mask_w1[77]
  PIN w_mask_w1[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.265 0.070 62.335 ;
    END
  END w_mask_w1[78]
  PIN w_mask_w1[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.685 0.070 62.755 ;
    END
  END w_mask_w1[79]
  PIN w_mask_w1[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.105 0.070 63.175 ;
    END
  END w_mask_w1[80]
  PIN w_mask_w1[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.525 0.070 63.595 ;
    END
  END w_mask_w1[81]
  PIN w_mask_w1[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.945 0.070 64.015 ;
    END
  END w_mask_w1[82]
  PIN w_mask_w1[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.365 0.070 64.435 ;
    END
  END w_mask_w1[83]
  PIN w_mask_w1[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.785 0.070 64.855 ;
    END
  END w_mask_w1[84]
  PIN w_mask_w1[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.205 0.070 65.275 ;
    END
  END w_mask_w1[85]
  PIN w_mask_w1[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.625 0.070 65.695 ;
    END
  END w_mask_w1[86]
  PIN w_mask_w1[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.045 0.070 66.115 ;
    END
  END w_mask_w1[87]
  PIN w_mask_w1[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.465 0.070 66.535 ;
    END
  END w_mask_w1[88]
  PIN w_mask_w1[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.885 0.070 66.955 ;
    END
  END w_mask_w1[89]
  PIN w_mask_w1[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.305 0.070 67.375 ;
    END
  END w_mask_w1[90]
  PIN w_mask_w1[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.725 0.070 67.795 ;
    END
  END w_mask_w1[91]
  PIN w_mask_w1[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.145 0.070 68.215 ;
    END
  END w_mask_w1[92]
  PIN w_mask_w1[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.565 0.070 68.635 ;
    END
  END w_mask_w1[93]
  PIN w_mask_w1[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.985 0.070 69.055 ;
    END
  END w_mask_w1[94]
  PIN w_mask_w1[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.405 0.070 69.475 ;
    END
  END w_mask_w1[95]
  PIN w_mask_w1[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.825 0.070 69.895 ;
    END
  END w_mask_w1[96]
  PIN w_mask_w1[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.245 0.070 70.315 ;
    END
  END w_mask_w1[97]
  PIN w_mask_w1[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.665 0.070 70.735 ;
    END
  END w_mask_w1[98]
  PIN w_mask_w1[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.085 0.070 71.155 ;
    END
  END w_mask_w1[99]
  PIN w_mask_w1[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.505 0.070 71.575 ;
    END
  END w_mask_w1[100]
  PIN w_mask_w1[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.925 0.070 71.995 ;
    END
  END w_mask_w1[101]
  PIN w_mask_w1[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.345 0.070 72.415 ;
    END
  END w_mask_w1[102]
  PIN w_mask_w1[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.765 0.070 72.835 ;
    END
  END w_mask_w1[103]
  PIN w_mask_w1[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.185 0.070 73.255 ;
    END
  END w_mask_w1[104]
  PIN w_mask_w1[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.605 0.070 73.675 ;
    END
  END w_mask_w1[105]
  PIN w_mask_w1[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.025 0.070 74.095 ;
    END
  END w_mask_w1[106]
  PIN w_mask_w1[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.445 0.070 74.515 ;
    END
  END w_mask_w1[107]
  PIN w_mask_w1[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.865 0.070 74.935 ;
    END
  END w_mask_w1[108]
  PIN w_mask_w1[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.285 0.070 75.355 ;
    END
  END w_mask_w1[109]
  PIN w_mask_w1[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.705 0.070 75.775 ;
    END
  END w_mask_w1[110]
  PIN w_mask_w1[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.125 0.070 76.195 ;
    END
  END w_mask_w1[111]
  PIN w_mask_w1[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.545 0.070 76.615 ;
    END
  END w_mask_w1[112]
  PIN w_mask_w1[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.965 0.070 77.035 ;
    END
  END w_mask_w1[113]
  PIN w_mask_w1[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.385 0.070 77.455 ;
    END
  END w_mask_w1[114]
  PIN w_mask_w1[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END w_mask_w1[115]
  PIN w_mask_w1[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.225 0.070 78.295 ;
    END
  END w_mask_w1[116]
  PIN w_mask_w1[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.645 0.070 78.715 ;
    END
  END w_mask_w1[117]
  PIN w_mask_w1[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.065 0.070 79.135 ;
    END
  END w_mask_w1[118]
  PIN w_mask_w1[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.485 0.070 79.555 ;
    END
  END w_mask_w1[119]
  PIN w_mask_w1[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.905 0.070 79.975 ;
    END
  END w_mask_w1[120]
  PIN w_mask_w1[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.325 0.070 80.395 ;
    END
  END w_mask_w1[121]
  PIN w_mask_w1[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.745 0.070 80.815 ;
    END
  END w_mask_w1[122]
  PIN w_mask_w1[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.165 0.070 81.235 ;
    END
  END w_mask_w1[123]
  PIN w_mask_w1[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.585 0.070 81.655 ;
    END
  END w_mask_w1[124]
  PIN w_mask_w1[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.005 0.070 82.075 ;
    END
  END w_mask_w1[125]
  PIN w_mask_w1[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.425 0.070 82.495 ;
    END
  END w_mask_w1[126]
  PIN w_mask_w1[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.845 0.070 82.915 ;
    END
  END w_mask_w1[127]
  PIN w_mask_w1[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.265 0.070 83.335 ;
    END
  END w_mask_w1[128]
  PIN w_mask_w1[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.685 0.070 83.755 ;
    END
  END w_mask_w1[129]
  PIN w_mask_w1[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.105 0.070 84.175 ;
    END
  END w_mask_w1[130]
  PIN w_mask_w1[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.525 0.070 84.595 ;
    END
  END w_mask_w1[131]
  PIN w_mask_w1[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.945 0.070 85.015 ;
    END
  END w_mask_w1[132]
  PIN w_mask_w1[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.365 0.070 85.435 ;
    END
  END w_mask_w1[133]
  PIN w_mask_w1[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.785 0.070 85.855 ;
    END
  END w_mask_w1[134]
  PIN w_mask_w1[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.205 0.070 86.275 ;
    END
  END w_mask_w1[135]
  PIN w_mask_w1[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.625 0.070 86.695 ;
    END
  END w_mask_w1[136]
  PIN w_mask_w1[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.045 0.070 87.115 ;
    END
  END w_mask_w1[137]
  PIN w_mask_w1[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.465 0.070 87.535 ;
    END
  END w_mask_w1[138]
  PIN w_mask_w1[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.885 0.070 87.955 ;
    END
  END w_mask_w1[139]
  PIN w_mask_w1[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.305 0.070 88.375 ;
    END
  END w_mask_w1[140]
  PIN w_mask_w1[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.725 0.070 88.795 ;
    END
  END w_mask_w1[141]
  PIN w_mask_w1[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.145 0.070 89.215 ;
    END
  END w_mask_w1[142]
  PIN w_mask_w1[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.565 0.070 89.635 ;
    END
  END w_mask_w1[143]
  PIN w_mask_w1[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.985 0.070 90.055 ;
    END
  END w_mask_w1[144]
  PIN w_mask_w1[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.405 0.070 90.475 ;
    END
  END w_mask_w1[145]
  PIN w_mask_w1[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.825 0.070 90.895 ;
    END
  END w_mask_w1[146]
  PIN w_mask_w1[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.245 0.070 91.315 ;
    END
  END w_mask_w1[147]
  PIN w_mask_w1[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.665 0.070 91.735 ;
    END
  END w_mask_w1[148]
  PIN w_mask_w1[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.085 0.070 92.155 ;
    END
  END w_mask_w1[149]
  PIN w_mask_w1[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.505 0.070 92.575 ;
    END
  END w_mask_w1[150]
  PIN w_mask_w1[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.925 0.070 92.995 ;
    END
  END w_mask_w1[151]
  PIN w_mask_w1[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.345 0.070 93.415 ;
    END
  END w_mask_w1[152]
  PIN w_mask_w1[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.765 0.070 93.835 ;
    END
  END w_mask_w1[153]
  PIN w_mask_w1[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.185 0.070 94.255 ;
    END
  END w_mask_w1[154]
  PIN w_mask_w1[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.605 0.070 94.675 ;
    END
  END w_mask_w1[155]
  PIN w_mask_w1[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.025 0.070 95.095 ;
    END
  END w_mask_w1[156]
  PIN w_mask_w1[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.445 0.070 95.515 ;
    END
  END w_mask_w1[157]
  PIN w_mask_w1[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.865 0.070 95.935 ;
    END
  END w_mask_w1[158]
  PIN w_mask_w1[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.285 0.070 96.355 ;
    END
  END w_mask_w1[159]
  PIN w_mask_w1[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.705 0.070 96.775 ;
    END
  END w_mask_w1[160]
  PIN w_mask_w1[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.125 0.070 97.195 ;
    END
  END w_mask_w1[161]
  PIN w_mask_w1[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.545 0.070 97.615 ;
    END
  END w_mask_w1[162]
  PIN w_mask_w1[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.965 0.070 98.035 ;
    END
  END w_mask_w1[163]
  PIN w_mask_w1[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.385 0.070 98.455 ;
    END
  END w_mask_w1[164]
  PIN w_mask_w1[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.805 0.070 98.875 ;
    END
  END w_mask_w1[165]
  PIN w_mask_w1[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.225 0.070 99.295 ;
    END
  END w_mask_w1[166]
  PIN w_mask_w1[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.645 0.070 99.715 ;
    END
  END w_mask_w1[167]
  PIN w_mask_w1[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.065 0.070 100.135 ;
    END
  END w_mask_w1[168]
  PIN w_mask_w1[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.485 0.070 100.555 ;
    END
  END w_mask_w1[169]
  PIN w_mask_w1[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.905 0.070 100.975 ;
    END
  END w_mask_w1[170]
  PIN w_mask_w1[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.325 0.070 101.395 ;
    END
  END w_mask_w1[171]
  PIN w_mask_w1[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.745 0.070 101.815 ;
    END
  END w_mask_w1[172]
  PIN w_mask_w1[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.165 0.070 102.235 ;
    END
  END w_mask_w1[173]
  PIN w_mask_w1[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.585 0.070 102.655 ;
    END
  END w_mask_w1[174]
  PIN w_mask_w1[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.005 0.070 103.075 ;
    END
  END w_mask_w1[175]
  PIN w_mask_w1[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.425 0.070 103.495 ;
    END
  END w_mask_w1[176]
  PIN w_mask_w1[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.845 0.070 103.915 ;
    END
  END w_mask_w1[177]
  PIN w_mask_w1[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.265 0.070 104.335 ;
    END
  END w_mask_w1[178]
  PIN w_mask_w1[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.685 0.070 104.755 ;
    END
  END w_mask_w1[179]
  PIN w_mask_w1[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.105 0.070 105.175 ;
    END
  END w_mask_w1[180]
  PIN w_mask_w1[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.525 0.070 105.595 ;
    END
  END w_mask_w1[181]
  PIN w_mask_w1[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.945 0.070 106.015 ;
    END
  END w_mask_w1[182]
  PIN w_mask_w1[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.365 0.070 106.435 ;
    END
  END w_mask_w1[183]
  PIN w_mask_w1[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.785 0.070 106.855 ;
    END
  END w_mask_w1[184]
  PIN w_mask_w1[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.205 0.070 107.275 ;
    END
  END w_mask_w1[185]
  PIN w_mask_w1[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.625 0.070 107.695 ;
    END
  END w_mask_w1[186]
  PIN w_mask_w1[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.045 0.070 108.115 ;
    END
  END w_mask_w1[187]
  PIN w_mask_w1[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.465 0.070 108.535 ;
    END
  END w_mask_w1[188]
  PIN w_mask_w1[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.885 0.070 108.955 ;
    END
  END w_mask_w1[189]
  PIN w_mask_w1[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.305 0.070 109.375 ;
    END
  END w_mask_w1[190]
  PIN w_mask_w1[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.725 0.070 109.795 ;
    END
  END w_mask_w1[191]
  PIN w_mask_w1[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.145 0.070 110.215 ;
    END
  END w_mask_w1[192]
  PIN w_mask_w1[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.565 0.070 110.635 ;
    END
  END w_mask_w1[193]
  PIN w_mask_w1[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.985 0.070 111.055 ;
    END
  END w_mask_w1[194]
  PIN w_mask_w1[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.405 0.070 111.475 ;
    END
  END w_mask_w1[195]
  PIN w_mask_w1[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.825 0.070 111.895 ;
    END
  END w_mask_w1[196]
  PIN w_mask_w1[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.245 0.070 112.315 ;
    END
  END w_mask_w1[197]
  PIN w_mask_w1[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.665 0.070 112.735 ;
    END
  END w_mask_w1[198]
  PIN w_mask_w1[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.085 0.070 113.155 ;
    END
  END w_mask_w1[199]
  PIN w_mask_w1[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.505 0.070 113.575 ;
    END
  END w_mask_w1[200]
  PIN w_mask_w1[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.925 0.070 113.995 ;
    END
  END w_mask_w1[201]
  PIN w_mask_w1[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.345 0.070 114.415 ;
    END
  END w_mask_w1[202]
  PIN w_mask_w1[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.765 0.070 114.835 ;
    END
  END w_mask_w1[203]
  PIN w_mask_w1[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.185 0.070 115.255 ;
    END
  END w_mask_w1[204]
  PIN w_mask_w1[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.605 0.070 115.675 ;
    END
  END w_mask_w1[205]
  PIN w_mask_w1[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.025 0.070 116.095 ;
    END
  END w_mask_w1[206]
  PIN w_mask_w1[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.445 0.070 116.515 ;
    END
  END w_mask_w1[207]
  PIN w_mask_w1[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.865 0.070 116.935 ;
    END
  END w_mask_w1[208]
  PIN w_mask_w1[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.285 0.070 117.355 ;
    END
  END w_mask_w1[209]
  PIN w_mask_w1[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.705 0.070 117.775 ;
    END
  END w_mask_w1[210]
  PIN w_mask_w1[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.125 0.070 118.195 ;
    END
  END w_mask_w1[211]
  PIN w_mask_w1[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.545 0.070 118.615 ;
    END
  END w_mask_w1[212]
  PIN w_mask_w1[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.965 0.070 119.035 ;
    END
  END w_mask_w1[213]
  PIN w_mask_w1[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.385 0.070 119.455 ;
    END
  END w_mask_w1[214]
  PIN w_mask_w1[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.805 0.070 119.875 ;
    END
  END w_mask_w1[215]
  PIN w_mask_w1[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.225 0.070 120.295 ;
    END
  END w_mask_w1[216]
  PIN w_mask_w1[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.645 0.070 120.715 ;
    END
  END w_mask_w1[217]
  PIN w_mask_w1[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.065 0.070 121.135 ;
    END
  END w_mask_w1[218]
  PIN w_mask_w1[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.485 0.070 121.555 ;
    END
  END w_mask_w1[219]
  PIN w_mask_w1[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.905 0.070 121.975 ;
    END
  END w_mask_w1[220]
  PIN w_mask_w1[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.325 0.070 122.395 ;
    END
  END w_mask_w1[221]
  PIN w_mask_w1[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.745 0.070 122.815 ;
    END
  END w_mask_w1[222]
  PIN w_mask_w1[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.165 0.070 123.235 ;
    END
  END w_mask_w1[223]
  PIN w_mask_w1[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.585 0.070 123.655 ;
    END
  END w_mask_w1[224]
  PIN w_mask_w1[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.005 0.070 124.075 ;
    END
  END w_mask_w1[225]
  PIN w_mask_w1[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.425 0.070 124.495 ;
    END
  END w_mask_w1[226]
  PIN w_mask_w1[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.845 0.070 124.915 ;
    END
  END w_mask_w1[227]
  PIN w_mask_w1[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.265 0.070 125.335 ;
    END
  END w_mask_w1[228]
  PIN w_mask_w1[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.685 0.070 125.755 ;
    END
  END w_mask_w1[229]
  PIN w_mask_w1[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.105 0.070 126.175 ;
    END
  END w_mask_w1[230]
  PIN w_mask_w1[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.525 0.070 126.595 ;
    END
  END w_mask_w1[231]
  PIN w_mask_w1[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.945 0.070 127.015 ;
    END
  END w_mask_w1[232]
  PIN w_mask_w1[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.365 0.070 127.435 ;
    END
  END w_mask_w1[233]
  PIN w_mask_w1[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.785 0.070 127.855 ;
    END
  END w_mask_w1[234]
  PIN w_mask_w1[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.205 0.070 128.275 ;
    END
  END w_mask_w1[235]
  PIN w_mask_w1[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.625 0.070 128.695 ;
    END
  END w_mask_w1[236]
  PIN w_mask_w1[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.045 0.070 129.115 ;
    END
  END w_mask_w1[237]
  PIN w_mask_w1[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.465 0.070 129.535 ;
    END
  END w_mask_w1[238]
  PIN w_mask_w1[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.885 0.070 129.955 ;
    END
  END w_mask_w1[239]
  PIN w_mask_w1[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.305 0.070 130.375 ;
    END
  END w_mask_w1[240]
  PIN w_mask_w1[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.725 0.070 130.795 ;
    END
  END w_mask_w1[241]
  PIN w_mask_w1[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.145 0.070 131.215 ;
    END
  END w_mask_w1[242]
  PIN w_mask_w1[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.565 0.070 131.635 ;
    END
  END w_mask_w1[243]
  PIN w_mask_w1[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.985 0.070 132.055 ;
    END
  END w_mask_w1[244]
  PIN w_mask_w1[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.405 0.070 132.475 ;
    END
  END w_mask_w1[245]
  PIN w_mask_w1[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.825 0.070 132.895 ;
    END
  END w_mask_w1[246]
  PIN w_mask_w1[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.245 0.070 133.315 ;
    END
  END w_mask_w1[247]
  PIN w_mask_w1[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.665 0.070 133.735 ;
    END
  END w_mask_w1[248]
  PIN w_mask_w1[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.085 0.070 134.155 ;
    END
  END w_mask_w1[249]
  PIN w_mask_w1[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.505 0.070 134.575 ;
    END
  END w_mask_w1[250]
  PIN w_mask_w1[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.925 0.070 134.995 ;
    END
  END w_mask_w1[251]
  PIN w_mask_w1[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.345 0.070 135.415 ;
    END
  END w_mask_w1[252]
  PIN w_mask_w1[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.765 0.070 135.835 ;
    END
  END w_mask_w1[253]
  PIN w_mask_w1[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.185 0.070 136.255 ;
    END
  END w_mask_w1[254]
  PIN w_mask_w1[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.605 0.070 136.675 ;
    END
  END w_mask_w1[255]
  PIN w_mask_w1[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.025 0.070 137.095 ;
    END
  END w_mask_w1[256]
  PIN w_mask_w1[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.445 0.070 137.515 ;
    END
  END w_mask_w1[257]
  PIN w_mask_w1[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.865 0.070 137.935 ;
    END
  END w_mask_w1[258]
  PIN w_mask_w1[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.285 0.070 138.355 ;
    END
  END w_mask_w1[259]
  PIN w_mask_w1[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.705 0.070 138.775 ;
    END
  END w_mask_w1[260]
  PIN w_mask_w1[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.125 0.070 139.195 ;
    END
  END w_mask_w1[261]
  PIN w_mask_w1[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.545 0.070 139.615 ;
    END
  END w_mask_w1[262]
  PIN w_mask_w1[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.965 0.070 140.035 ;
    END
  END w_mask_w1[263]
  PIN w_mask_w1[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.385 0.070 140.455 ;
    END
  END w_mask_w1[264]
  PIN w_mask_w1[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.805 0.070 140.875 ;
    END
  END w_mask_w1[265]
  PIN w_mask_w1[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.225 0.070 141.295 ;
    END
  END w_mask_w1[266]
  PIN w_mask_w1[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.645 0.070 141.715 ;
    END
  END w_mask_w1[267]
  PIN w_mask_w1[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.065 0.070 142.135 ;
    END
  END w_mask_w1[268]
  PIN w_mask_w1[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.485 0.070 142.555 ;
    END
  END w_mask_w1[269]
  PIN w_mask_w1[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.905 0.070 142.975 ;
    END
  END w_mask_w1[270]
  PIN w_mask_w1[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.325 0.070 143.395 ;
    END
  END w_mask_w1[271]
  PIN w_mask_w1[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.745 0.070 143.815 ;
    END
  END w_mask_w1[272]
  PIN w_mask_w1[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.165 0.070 144.235 ;
    END
  END w_mask_w1[273]
  PIN w_mask_w1[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.585 0.070 144.655 ;
    END
  END w_mask_w1[274]
  PIN w_mask_w1[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.005 0.070 145.075 ;
    END
  END w_mask_w1[275]
  PIN w_mask_w1[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.425 0.070 145.495 ;
    END
  END w_mask_w1[276]
  PIN w_mask_w1[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.845 0.070 145.915 ;
    END
  END w_mask_w1[277]
  PIN w_mask_w1[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.265 0.070 146.335 ;
    END
  END w_mask_w1[278]
  PIN w_mask_w1[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.685 0.070 146.755 ;
    END
  END w_mask_w1[279]
  PIN w_mask_w1[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.105 0.070 147.175 ;
    END
  END w_mask_w1[280]
  PIN w_mask_w1[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.525 0.070 147.595 ;
    END
  END w_mask_w1[281]
  PIN w_mask_w1[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.945 0.070 148.015 ;
    END
  END w_mask_w1[282]
  PIN w_mask_w1[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.365 0.070 148.435 ;
    END
  END w_mask_w1[283]
  PIN w_mask_w1[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.785 0.070 148.855 ;
    END
  END w_mask_w1[284]
  PIN w_mask_w1[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.205 0.070 149.275 ;
    END
  END w_mask_w1[285]
  PIN w_mask_w1[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.625 0.070 149.695 ;
    END
  END w_mask_w1[286]
  PIN w_mask_w1[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.045 0.070 150.115 ;
    END
  END w_mask_w1[287]
  PIN w_mask_w1[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.465 0.070 150.535 ;
    END
  END w_mask_w1[288]
  PIN w_mask_w1[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.885 0.070 150.955 ;
    END
  END w_mask_w1[289]
  PIN w_mask_w1[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.305 0.070 151.375 ;
    END
  END w_mask_w1[290]
  PIN w_mask_w1[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.725 0.070 151.795 ;
    END
  END w_mask_w1[291]
  PIN w_mask_w1[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.145 0.070 152.215 ;
    END
  END w_mask_w1[292]
  PIN w_mask_w1[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.565 0.070 152.635 ;
    END
  END w_mask_w1[293]
  PIN w_mask_w1[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.985 0.070 153.055 ;
    END
  END w_mask_w1[294]
  PIN w_mask_w1[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.405 0.070 153.475 ;
    END
  END w_mask_w1[295]
  PIN w_mask_w1[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.825 0.070 153.895 ;
    END
  END w_mask_w1[296]
  PIN w_mask_w1[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.245 0.070 154.315 ;
    END
  END w_mask_w1[297]
  PIN w_mask_w1[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.665 0.070 154.735 ;
    END
  END w_mask_w1[298]
  PIN w_mask_w1[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.085 0.070 155.155 ;
    END
  END w_mask_w1[299]
  PIN w_mask_w1[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.505 0.070 155.575 ;
    END
  END w_mask_w1[300]
  PIN w_mask_w1[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.925 0.070 155.995 ;
    END
  END w_mask_w1[301]
  PIN w_mask_w1[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.345 0.070 156.415 ;
    END
  END w_mask_w1[302]
  PIN w_mask_w1[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.765 0.070 156.835 ;
    END
  END w_mask_w1[303]
  PIN w_mask_w1[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.185 0.070 157.255 ;
    END
  END w_mask_w1[304]
  PIN w_mask_w1[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.605 0.070 157.675 ;
    END
  END w_mask_w1[305]
  PIN w_mask_w1[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.025 0.070 158.095 ;
    END
  END w_mask_w1[306]
  PIN w_mask_w1[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.445 0.070 158.515 ;
    END
  END w_mask_w1[307]
  PIN w_mask_w1[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.865 0.070 158.935 ;
    END
  END w_mask_w1[308]
  PIN w_mask_w1[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.285 0.070 159.355 ;
    END
  END w_mask_w1[309]
  PIN w_mask_w1[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.705 0.070 159.775 ;
    END
  END w_mask_w1[310]
  PIN w_mask_w1[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.125 0.070 160.195 ;
    END
  END w_mask_w1[311]
  PIN w_mask_w1[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.545 0.070 160.615 ;
    END
  END w_mask_w1[312]
  PIN w_mask_w1[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.965 0.070 161.035 ;
    END
  END w_mask_w1[313]
  PIN w_mask_w1[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.385 0.070 161.455 ;
    END
  END w_mask_w1[314]
  PIN w_mask_w1[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.805 0.070 161.875 ;
    END
  END w_mask_w1[315]
  PIN w_mask_w1[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.225 0.070 162.295 ;
    END
  END w_mask_w1[316]
  PIN w_mask_w1[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.645 0.070 162.715 ;
    END
  END w_mask_w1[317]
  PIN w_mask_w1[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.065 0.070 163.135 ;
    END
  END w_mask_w1[318]
  PIN w_mask_w1[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.485 0.070 163.555 ;
    END
  END w_mask_w1[319]
  PIN w_mask_w1[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.905 0.070 163.975 ;
    END
  END w_mask_w1[320]
  PIN w_mask_w1[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.325 0.070 164.395 ;
    END
  END w_mask_w1[321]
  PIN w_mask_w1[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.745 0.070 164.815 ;
    END
  END w_mask_w1[322]
  PIN w_mask_w1[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.165 0.070 165.235 ;
    END
  END w_mask_w1[323]
  PIN w_mask_w1[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.585 0.070 165.655 ;
    END
  END w_mask_w1[324]
  PIN w_mask_w1[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.005 0.070 166.075 ;
    END
  END w_mask_w1[325]
  PIN w_mask_w1[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.425 0.070 166.495 ;
    END
  END w_mask_w1[326]
  PIN w_mask_w1[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.845 0.070 166.915 ;
    END
  END w_mask_w1[327]
  PIN w_mask_w1[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.265 0.070 167.335 ;
    END
  END w_mask_w1[328]
  PIN w_mask_w1[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.685 0.070 167.755 ;
    END
  END w_mask_w1[329]
  PIN w_mask_w1[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.105 0.070 168.175 ;
    END
  END w_mask_w1[330]
  PIN w_mask_w1[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.525 0.070 168.595 ;
    END
  END w_mask_w1[331]
  PIN w_mask_w1[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.945 0.070 169.015 ;
    END
  END w_mask_w1[332]
  PIN w_mask_w1[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.365 0.070 169.435 ;
    END
  END w_mask_w1[333]
  PIN w_mask_w1[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.785 0.070 169.855 ;
    END
  END w_mask_w1[334]
  PIN w_mask_w1[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.205 0.070 170.275 ;
    END
  END w_mask_w1[335]
  PIN w_mask_w1[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.625 0.070 170.695 ;
    END
  END w_mask_w1[336]
  PIN w_mask_w1[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.045 0.070 171.115 ;
    END
  END w_mask_w1[337]
  PIN w_mask_w1[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.465 0.070 171.535 ;
    END
  END w_mask_w1[338]
  PIN w_mask_w1[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.885 0.070 171.955 ;
    END
  END w_mask_w1[339]
  PIN w_mask_w1[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.305 0.070 172.375 ;
    END
  END w_mask_w1[340]
  PIN w_mask_w1[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.725 0.070 172.795 ;
    END
  END w_mask_w1[341]
  PIN w_mask_w1[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.145 0.070 173.215 ;
    END
  END w_mask_w1[342]
  PIN w_mask_w1[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.565 0.070 173.635 ;
    END
  END w_mask_w1[343]
  PIN w_mask_w1[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.985 0.070 174.055 ;
    END
  END w_mask_w1[344]
  PIN w_mask_w1[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.405 0.070 174.475 ;
    END
  END w_mask_w1[345]
  PIN w_mask_w1[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.825 0.070 174.895 ;
    END
  END w_mask_w1[346]
  PIN w_mask_w1[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.245 0.070 175.315 ;
    END
  END w_mask_w1[347]
  PIN w_mask_w1[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.665 0.070 175.735 ;
    END
  END w_mask_w1[348]
  PIN w_mask_w1[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.085 0.070 176.155 ;
    END
  END w_mask_w1[349]
  PIN w_mask_w1[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.505 0.070 176.575 ;
    END
  END w_mask_w1[350]
  PIN w_mask_w1[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.925 0.070 176.995 ;
    END
  END w_mask_w1[351]
  PIN w_mask_w1[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.345 0.070 177.415 ;
    END
  END w_mask_w1[352]
  PIN w_mask_w1[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.765 0.070 177.835 ;
    END
  END w_mask_w1[353]
  PIN w_mask_w1[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.185 0.070 178.255 ;
    END
  END w_mask_w1[354]
  PIN w_mask_w1[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.605 0.070 178.675 ;
    END
  END w_mask_w1[355]
  PIN w_mask_w1[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.025 0.070 179.095 ;
    END
  END w_mask_w1[356]
  PIN w_mask_w1[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.445 0.070 179.515 ;
    END
  END w_mask_w1[357]
  PIN w_mask_w1[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.865 0.070 179.935 ;
    END
  END w_mask_w1[358]
  PIN w_mask_w1[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.285 0.070 180.355 ;
    END
  END w_mask_w1[359]
  PIN w_mask_w1[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.705 0.070 180.775 ;
    END
  END w_mask_w1[360]
  PIN w_mask_w1[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.125 0.070 181.195 ;
    END
  END w_mask_w1[361]
  PIN w_mask_w1[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.545 0.070 181.615 ;
    END
  END w_mask_w1[362]
  PIN w_mask_w1[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.965 0.070 182.035 ;
    END
  END w_mask_w1[363]
  PIN w_mask_w1[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.385 0.070 182.455 ;
    END
  END w_mask_w1[364]
  PIN w_mask_w1[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.805 0.070 182.875 ;
    END
  END w_mask_w1[365]
  PIN w_mask_w1[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.225 0.070 183.295 ;
    END
  END w_mask_w1[366]
  PIN w_mask_w1[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.645 0.070 183.715 ;
    END
  END w_mask_w1[367]
  PIN w_mask_w1[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.065 0.070 184.135 ;
    END
  END w_mask_w1[368]
  PIN w_mask_w1[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.485 0.070 184.555 ;
    END
  END w_mask_w1[369]
  PIN w_mask_w1[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.905 0.070 184.975 ;
    END
  END w_mask_w1[370]
  PIN w_mask_w1[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.325 0.070 185.395 ;
    END
  END w_mask_w1[371]
  PIN w_mask_w1[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.745 0.070 185.815 ;
    END
  END w_mask_w1[372]
  PIN w_mask_w1[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.165 0.070 186.235 ;
    END
  END w_mask_w1[373]
  PIN w_mask_w1[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.585 0.070 186.655 ;
    END
  END w_mask_w1[374]
  PIN w_mask_w1[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.005 0.070 187.075 ;
    END
  END w_mask_w1[375]
  PIN w_mask_w1[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.425 0.070 187.495 ;
    END
  END w_mask_w1[376]
  PIN w_mask_w1[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.845 0.070 187.915 ;
    END
  END w_mask_w1[377]
  PIN w_mask_w1[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.265 0.070 188.335 ;
    END
  END w_mask_w1[378]
  PIN w_mask_w1[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.685 0.070 188.755 ;
    END
  END w_mask_w1[379]
  PIN w_mask_w1[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.105 0.070 189.175 ;
    END
  END w_mask_w1[380]
  PIN w_mask_w1[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.525 0.070 189.595 ;
    END
  END w_mask_w1[381]
  PIN w_mask_w1[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.945 0.070 190.015 ;
    END
  END w_mask_w1[382]
  PIN w_mask_w1[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.365 0.070 190.435 ;
    END
  END w_mask_w1[383]
  PIN w_mask_w1[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.785 0.070 190.855 ;
    END
  END w_mask_w1[384]
  PIN w_mask_w1[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.205 0.070 191.275 ;
    END
  END w_mask_w1[385]
  PIN w_mask_w1[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.625 0.070 191.695 ;
    END
  END w_mask_w1[386]
  PIN w_mask_w1[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.045 0.070 192.115 ;
    END
  END w_mask_w1[387]
  PIN w_mask_w1[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.465 0.070 192.535 ;
    END
  END w_mask_w1[388]
  PIN w_mask_w1[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.885 0.070 192.955 ;
    END
  END w_mask_w1[389]
  PIN w_mask_w1[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.305 0.070 193.375 ;
    END
  END w_mask_w1[390]
  PIN w_mask_w1[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.725 0.070 193.795 ;
    END
  END w_mask_w1[391]
  PIN w_mask_w1[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.145 0.070 194.215 ;
    END
  END w_mask_w1[392]
  PIN w_mask_w1[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.565 0.070 194.635 ;
    END
  END w_mask_w1[393]
  PIN w_mask_w1[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.985 0.070 195.055 ;
    END
  END w_mask_w1[394]
  PIN w_mask_w1[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.405 0.070 195.475 ;
    END
  END w_mask_w1[395]
  PIN w_mask_w1[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.825 0.070 195.895 ;
    END
  END w_mask_w1[396]
  PIN w_mask_w1[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.245 0.070 196.315 ;
    END
  END w_mask_w1[397]
  PIN w_mask_w1[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.665 0.070 196.735 ;
    END
  END w_mask_w1[398]
  PIN w_mask_w1[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.085 0.070 197.155 ;
    END
  END w_mask_w1[399]
  PIN w_mask_w1[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.505 0.070 197.575 ;
    END
  END w_mask_w1[400]
  PIN w_mask_w1[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.925 0.070 197.995 ;
    END
  END w_mask_w1[401]
  PIN w_mask_w1[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.345 0.070 198.415 ;
    END
  END w_mask_w1[402]
  PIN w_mask_w1[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.765 0.070 198.835 ;
    END
  END w_mask_w1[403]
  PIN w_mask_w1[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.185 0.070 199.255 ;
    END
  END w_mask_w1[404]
  PIN w_mask_w1[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.605 0.070 199.675 ;
    END
  END w_mask_w1[405]
  PIN w_mask_w1[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.025 0.070 200.095 ;
    END
  END w_mask_w1[406]
  PIN w_mask_w1[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.445 0.070 200.515 ;
    END
  END w_mask_w1[407]
  PIN w_mask_w1[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.865 0.070 200.935 ;
    END
  END w_mask_w1[408]
  PIN w_mask_w1[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.285 0.070 201.355 ;
    END
  END w_mask_w1[409]
  PIN w_mask_w1[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.705 0.070 201.775 ;
    END
  END w_mask_w1[410]
  PIN w_mask_w1[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.125 0.070 202.195 ;
    END
  END w_mask_w1[411]
  PIN w_mask_w1[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.545 0.070 202.615 ;
    END
  END w_mask_w1[412]
  PIN w_mask_w1[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.965 0.070 203.035 ;
    END
  END w_mask_w1[413]
  PIN w_mask_w1[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.385 0.070 203.455 ;
    END
  END w_mask_w1[414]
  PIN w_mask_w1[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.805 0.070 203.875 ;
    END
  END w_mask_w1[415]
  PIN w_mask_w1[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.225 0.070 204.295 ;
    END
  END w_mask_w1[416]
  PIN w_mask_w1[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.645 0.070 204.715 ;
    END
  END w_mask_w1[417]
  PIN w_mask_w1[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.065 0.070 205.135 ;
    END
  END w_mask_w1[418]
  PIN w_mask_w1[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.485 0.070 205.555 ;
    END
  END w_mask_w1[419]
  PIN w_mask_w1[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.905 0.070 205.975 ;
    END
  END w_mask_w1[420]
  PIN w_mask_w1[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.325 0.070 206.395 ;
    END
  END w_mask_w1[421]
  PIN w_mask_w1[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.745 0.070 206.815 ;
    END
  END w_mask_w1[422]
  PIN w_mask_w1[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.165 0.070 207.235 ;
    END
  END w_mask_w1[423]
  PIN w_mask_w1[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.585 0.070 207.655 ;
    END
  END w_mask_w1[424]
  PIN w_mask_w1[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.005 0.070 208.075 ;
    END
  END w_mask_w1[425]
  PIN w_mask_w1[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.425 0.070 208.495 ;
    END
  END w_mask_w1[426]
  PIN w_mask_w1[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.845 0.070 208.915 ;
    END
  END w_mask_w1[427]
  PIN w_mask_w1[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.265 0.070 209.335 ;
    END
  END w_mask_w1[428]
  PIN w_mask_w1[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.685 0.070 209.755 ;
    END
  END w_mask_w1[429]
  PIN w_mask_w1[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.105 0.070 210.175 ;
    END
  END w_mask_w1[430]
  PIN w_mask_w1[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.525 0.070 210.595 ;
    END
  END w_mask_w1[431]
  PIN w_mask_w1[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.945 0.070 211.015 ;
    END
  END w_mask_w1[432]
  PIN w_mask_w1[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.365 0.070 211.435 ;
    END
  END w_mask_w1[433]
  PIN w_mask_w1[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.785 0.070 211.855 ;
    END
  END w_mask_w1[434]
  PIN w_mask_w1[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.205 0.070 212.275 ;
    END
  END w_mask_w1[435]
  PIN w_mask_w1[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.625 0.070 212.695 ;
    END
  END w_mask_w1[436]
  PIN w_mask_w1[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.045 0.070 213.115 ;
    END
  END w_mask_w1[437]
  PIN w_mask_w1[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.465 0.070 213.535 ;
    END
  END w_mask_w1[438]
  PIN w_mask_w1[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.885 0.070 213.955 ;
    END
  END w_mask_w1[439]
  PIN w_mask_w1[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.305 0.070 214.375 ;
    END
  END w_mask_w1[440]
  PIN w_mask_w1[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.725 0.070 214.795 ;
    END
  END w_mask_w1[441]
  PIN w_mask_w1[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.145 0.070 215.215 ;
    END
  END w_mask_w1[442]
  PIN w_mask_w1[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.565 0.070 215.635 ;
    END
  END w_mask_w1[443]
  PIN w_mask_w1[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.985 0.070 216.055 ;
    END
  END w_mask_w1[444]
  PIN w_mask_w1[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.405 0.070 216.475 ;
    END
  END w_mask_w1[445]
  PIN w_mask_w1[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.825 0.070 216.895 ;
    END
  END w_mask_w1[446]
  PIN w_mask_w1[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.245 0.070 217.315 ;
    END
  END w_mask_w1[447]
  PIN w_mask_w1[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.665 0.070 217.735 ;
    END
  END w_mask_w1[448]
  PIN w_mask_w1[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.085 0.070 218.155 ;
    END
  END w_mask_w1[449]
  PIN w_mask_w1[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.505 0.070 218.575 ;
    END
  END w_mask_w1[450]
  PIN w_mask_w1[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.925 0.070 218.995 ;
    END
  END w_mask_w1[451]
  PIN w_mask_w1[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.345 0.070 219.415 ;
    END
  END w_mask_w1[452]
  PIN w_mask_w1[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.765 0.070 219.835 ;
    END
  END w_mask_w1[453]
  PIN w_mask_w1[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.185 0.070 220.255 ;
    END
  END w_mask_w1[454]
  PIN w_mask_w1[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.605 0.070 220.675 ;
    END
  END w_mask_w1[455]
  PIN w_mask_w1[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.025 0.070 221.095 ;
    END
  END w_mask_w1[456]
  PIN w_mask_w1[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.445 0.070 221.515 ;
    END
  END w_mask_w1[457]
  PIN w_mask_w1[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.865 0.070 221.935 ;
    END
  END w_mask_w1[458]
  PIN w_mask_w1[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.285 0.070 222.355 ;
    END
  END w_mask_w1[459]
  PIN w_mask_w1[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.705 0.070 222.775 ;
    END
  END w_mask_w1[460]
  PIN w_mask_w1[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.125 0.070 223.195 ;
    END
  END w_mask_w1[461]
  PIN w_mask_w1[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.545 0.070 223.615 ;
    END
  END w_mask_w1[462]
  PIN w_mask_w1[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.965 0.070 224.035 ;
    END
  END w_mask_w1[463]
  PIN w_mask_w1[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.385 0.070 224.455 ;
    END
  END w_mask_w1[464]
  PIN w_mask_w1[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.805 0.070 224.875 ;
    END
  END w_mask_w1[465]
  PIN w_mask_w1[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.225 0.070 225.295 ;
    END
  END w_mask_w1[466]
  PIN w_mask_w1[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.645 0.070 225.715 ;
    END
  END w_mask_w1[467]
  PIN w_mask_w1[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.065 0.070 226.135 ;
    END
  END w_mask_w1[468]
  PIN w_mask_w1[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.485 0.070 226.555 ;
    END
  END w_mask_w1[469]
  PIN w_mask_w1[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.905 0.070 226.975 ;
    END
  END w_mask_w1[470]
  PIN w_mask_w1[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.325 0.070 227.395 ;
    END
  END w_mask_w1[471]
  PIN w_mask_w1[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.745 0.070 227.815 ;
    END
  END w_mask_w1[472]
  PIN w_mask_w1[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.165 0.070 228.235 ;
    END
  END w_mask_w1[473]
  PIN w_mask_w1[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.585 0.070 228.655 ;
    END
  END w_mask_w1[474]
  PIN w_mask_w1[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.005 0.070 229.075 ;
    END
  END w_mask_w1[475]
  PIN w_mask_w1[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.425 0.070 229.495 ;
    END
  END w_mask_w1[476]
  PIN w_mask_w1[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.845 0.070 229.915 ;
    END
  END w_mask_w1[477]
  PIN w_mask_w1[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.265 0.070 230.335 ;
    END
  END w_mask_w1[478]
  PIN w_mask_w1[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.685 0.070 230.755 ;
    END
  END w_mask_w1[479]
  PIN w_mask_w1[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.105 0.070 231.175 ;
    END
  END w_mask_w1[480]
  PIN w_mask_w1[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.525 0.070 231.595 ;
    END
  END w_mask_w1[481]
  PIN w_mask_w1[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.945 0.070 232.015 ;
    END
  END w_mask_w1[482]
  PIN w_mask_w1[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.365 0.070 232.435 ;
    END
  END w_mask_w1[483]
  PIN w_mask_w1[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.785 0.070 232.855 ;
    END
  END w_mask_w1[484]
  PIN w_mask_w1[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.205 0.070 233.275 ;
    END
  END w_mask_w1[485]
  PIN w_mask_w1[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.625 0.070 233.695 ;
    END
  END w_mask_w1[486]
  PIN w_mask_w1[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.045 0.070 234.115 ;
    END
  END w_mask_w1[487]
  PIN w_mask_w1[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.465 0.070 234.535 ;
    END
  END w_mask_w1[488]
  PIN w_mask_w1[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.885 0.070 234.955 ;
    END
  END w_mask_w1[489]
  PIN w_mask_w1[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.305 0.070 235.375 ;
    END
  END w_mask_w1[490]
  PIN w_mask_w1[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.725 0.070 235.795 ;
    END
  END w_mask_w1[491]
  PIN w_mask_w1[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.145 0.070 236.215 ;
    END
  END w_mask_w1[492]
  PIN w_mask_w1[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.565 0.070 236.635 ;
    END
  END w_mask_w1[493]
  PIN w_mask_w1[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.985 0.070 237.055 ;
    END
  END w_mask_w1[494]
  PIN w_mask_w1[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.405 0.070 237.475 ;
    END
  END w_mask_w1[495]
  PIN w_mask_w1[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.825 0.070 237.895 ;
    END
  END w_mask_w1[496]
  PIN w_mask_w1[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.245 0.070 238.315 ;
    END
  END w_mask_w1[497]
  PIN w_mask_w1[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.665 0.070 238.735 ;
    END
  END w_mask_w1[498]
  PIN w_mask_w1[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.085 0.070 239.155 ;
    END
  END w_mask_w1[499]
  PIN w_mask_w1[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.505 0.070 239.575 ;
    END
  END w_mask_w1[500]
  PIN w_mask_w1[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.925 0.070 239.995 ;
    END
  END w_mask_w1[501]
  PIN w_mask_w1[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.345 0.070 240.415 ;
    END
  END w_mask_w1[502]
  PIN w_mask_w1[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.765 0.070 240.835 ;
    END
  END w_mask_w1[503]
  PIN w_mask_w1[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.185 0.070 241.255 ;
    END
  END w_mask_w1[504]
  PIN w_mask_w1[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.605 0.070 241.675 ;
    END
  END w_mask_w1[505]
  PIN w_mask_w1[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.025 0.070 242.095 ;
    END
  END w_mask_w1[506]
  PIN w_mask_w1[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.445 0.070 242.515 ;
    END
  END w_mask_w1[507]
  PIN w_mask_w1[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.865 0.070 242.935 ;
    END
  END w_mask_w1[508]
  PIN w_mask_w1[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.285 0.070 243.355 ;
    END
  END w_mask_w1[509]
  PIN w_mask_w1[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.705 0.070 243.775 ;
    END
  END w_mask_w1[510]
  PIN w_mask_w1[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.125 0.070 244.195 ;
    END
  END w_mask_w1[511]
  PIN rd_out_r1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.685 0.070 272.755 ;
    END
  END rd_out_r1[0]
  PIN rd_out_r1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.105 0.070 273.175 ;
    END
  END rd_out_r1[1]
  PIN rd_out_r1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.525 0.070 273.595 ;
    END
  END rd_out_r1[2]
  PIN rd_out_r1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.945 0.070 274.015 ;
    END
  END rd_out_r1[3]
  PIN rd_out_r1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.365 0.070 274.435 ;
    END
  END rd_out_r1[4]
  PIN rd_out_r1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.785 0.070 274.855 ;
    END
  END rd_out_r1[5]
  PIN rd_out_r1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.205 0.070 275.275 ;
    END
  END rd_out_r1[6]
  PIN rd_out_r1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.625 0.070 275.695 ;
    END
  END rd_out_r1[7]
  PIN rd_out_r1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.045 0.070 276.115 ;
    END
  END rd_out_r1[8]
  PIN rd_out_r1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.465 0.070 276.535 ;
    END
  END rd_out_r1[9]
  PIN rd_out_r1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.885 0.070 276.955 ;
    END
  END rd_out_r1[10]
  PIN rd_out_r1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.305 0.070 277.375 ;
    END
  END rd_out_r1[11]
  PIN rd_out_r1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.725 0.070 277.795 ;
    END
  END rd_out_r1[12]
  PIN rd_out_r1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.145 0.070 278.215 ;
    END
  END rd_out_r1[13]
  PIN rd_out_r1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.565 0.070 278.635 ;
    END
  END rd_out_r1[14]
  PIN rd_out_r1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.985 0.070 279.055 ;
    END
  END rd_out_r1[15]
  PIN rd_out_r1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.405 0.070 279.475 ;
    END
  END rd_out_r1[16]
  PIN rd_out_r1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.825 0.070 279.895 ;
    END
  END rd_out_r1[17]
  PIN rd_out_r1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.245 0.070 280.315 ;
    END
  END rd_out_r1[18]
  PIN rd_out_r1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.665 0.070 280.735 ;
    END
  END rd_out_r1[19]
  PIN rd_out_r1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.085 0.070 281.155 ;
    END
  END rd_out_r1[20]
  PIN rd_out_r1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.505 0.070 281.575 ;
    END
  END rd_out_r1[21]
  PIN rd_out_r1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.925 0.070 281.995 ;
    END
  END rd_out_r1[22]
  PIN rd_out_r1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.345 0.070 282.415 ;
    END
  END rd_out_r1[23]
  PIN rd_out_r1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.765 0.070 282.835 ;
    END
  END rd_out_r1[24]
  PIN rd_out_r1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.185 0.070 283.255 ;
    END
  END rd_out_r1[25]
  PIN rd_out_r1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.605 0.070 283.675 ;
    END
  END rd_out_r1[26]
  PIN rd_out_r1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.025 0.070 284.095 ;
    END
  END rd_out_r1[27]
  PIN rd_out_r1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.445 0.070 284.515 ;
    END
  END rd_out_r1[28]
  PIN rd_out_r1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.865 0.070 284.935 ;
    END
  END rd_out_r1[29]
  PIN rd_out_r1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.285 0.070 285.355 ;
    END
  END rd_out_r1[30]
  PIN rd_out_r1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.705 0.070 285.775 ;
    END
  END rd_out_r1[31]
  PIN rd_out_r1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.125 0.070 286.195 ;
    END
  END rd_out_r1[32]
  PIN rd_out_r1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.545 0.070 286.615 ;
    END
  END rd_out_r1[33]
  PIN rd_out_r1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.965 0.070 287.035 ;
    END
  END rd_out_r1[34]
  PIN rd_out_r1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.385 0.070 287.455 ;
    END
  END rd_out_r1[35]
  PIN rd_out_r1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.805 0.070 287.875 ;
    END
  END rd_out_r1[36]
  PIN rd_out_r1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.225 0.070 288.295 ;
    END
  END rd_out_r1[37]
  PIN rd_out_r1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.645 0.070 288.715 ;
    END
  END rd_out_r1[38]
  PIN rd_out_r1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.065 0.070 289.135 ;
    END
  END rd_out_r1[39]
  PIN rd_out_r1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.485 0.070 289.555 ;
    END
  END rd_out_r1[40]
  PIN rd_out_r1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.905 0.070 289.975 ;
    END
  END rd_out_r1[41]
  PIN rd_out_r1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.325 0.070 290.395 ;
    END
  END rd_out_r1[42]
  PIN rd_out_r1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.745 0.070 290.815 ;
    END
  END rd_out_r1[43]
  PIN rd_out_r1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.165 0.070 291.235 ;
    END
  END rd_out_r1[44]
  PIN rd_out_r1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.585 0.070 291.655 ;
    END
  END rd_out_r1[45]
  PIN rd_out_r1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.005 0.070 292.075 ;
    END
  END rd_out_r1[46]
  PIN rd_out_r1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.425 0.070 292.495 ;
    END
  END rd_out_r1[47]
  PIN rd_out_r1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.845 0.070 292.915 ;
    END
  END rd_out_r1[48]
  PIN rd_out_r1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.265 0.070 293.335 ;
    END
  END rd_out_r1[49]
  PIN rd_out_r1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.685 0.070 293.755 ;
    END
  END rd_out_r1[50]
  PIN rd_out_r1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.105 0.070 294.175 ;
    END
  END rd_out_r1[51]
  PIN rd_out_r1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.525 0.070 294.595 ;
    END
  END rd_out_r1[52]
  PIN rd_out_r1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.945 0.070 295.015 ;
    END
  END rd_out_r1[53]
  PIN rd_out_r1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.365 0.070 295.435 ;
    END
  END rd_out_r1[54]
  PIN rd_out_r1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.785 0.070 295.855 ;
    END
  END rd_out_r1[55]
  PIN rd_out_r1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.205 0.070 296.275 ;
    END
  END rd_out_r1[56]
  PIN rd_out_r1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.625 0.070 296.695 ;
    END
  END rd_out_r1[57]
  PIN rd_out_r1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.045 0.070 297.115 ;
    END
  END rd_out_r1[58]
  PIN rd_out_r1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.465 0.070 297.535 ;
    END
  END rd_out_r1[59]
  PIN rd_out_r1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.885 0.070 297.955 ;
    END
  END rd_out_r1[60]
  PIN rd_out_r1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.305 0.070 298.375 ;
    END
  END rd_out_r1[61]
  PIN rd_out_r1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.725 0.070 298.795 ;
    END
  END rd_out_r1[62]
  PIN rd_out_r1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.145 0.070 299.215 ;
    END
  END rd_out_r1[63]
  PIN rd_out_r1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.565 0.070 299.635 ;
    END
  END rd_out_r1[64]
  PIN rd_out_r1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.985 0.070 300.055 ;
    END
  END rd_out_r1[65]
  PIN rd_out_r1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.405 0.070 300.475 ;
    END
  END rd_out_r1[66]
  PIN rd_out_r1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.825 0.070 300.895 ;
    END
  END rd_out_r1[67]
  PIN rd_out_r1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.245 0.070 301.315 ;
    END
  END rd_out_r1[68]
  PIN rd_out_r1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.665 0.070 301.735 ;
    END
  END rd_out_r1[69]
  PIN rd_out_r1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.085 0.070 302.155 ;
    END
  END rd_out_r1[70]
  PIN rd_out_r1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.505 0.070 302.575 ;
    END
  END rd_out_r1[71]
  PIN rd_out_r1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.925 0.070 302.995 ;
    END
  END rd_out_r1[72]
  PIN rd_out_r1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.345 0.070 303.415 ;
    END
  END rd_out_r1[73]
  PIN rd_out_r1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.765 0.070 303.835 ;
    END
  END rd_out_r1[74]
  PIN rd_out_r1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.185 0.070 304.255 ;
    END
  END rd_out_r1[75]
  PIN rd_out_r1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.605 0.070 304.675 ;
    END
  END rd_out_r1[76]
  PIN rd_out_r1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.025 0.070 305.095 ;
    END
  END rd_out_r1[77]
  PIN rd_out_r1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.445 0.070 305.515 ;
    END
  END rd_out_r1[78]
  PIN rd_out_r1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.865 0.070 305.935 ;
    END
  END rd_out_r1[79]
  PIN rd_out_r1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.285 0.070 306.355 ;
    END
  END rd_out_r1[80]
  PIN rd_out_r1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.705 0.070 306.775 ;
    END
  END rd_out_r1[81]
  PIN rd_out_r1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.125 0.070 307.195 ;
    END
  END rd_out_r1[82]
  PIN rd_out_r1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.545 0.070 307.615 ;
    END
  END rd_out_r1[83]
  PIN rd_out_r1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.965 0.070 308.035 ;
    END
  END rd_out_r1[84]
  PIN rd_out_r1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.385 0.070 308.455 ;
    END
  END rd_out_r1[85]
  PIN rd_out_r1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.805 0.070 308.875 ;
    END
  END rd_out_r1[86]
  PIN rd_out_r1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.225 0.070 309.295 ;
    END
  END rd_out_r1[87]
  PIN rd_out_r1[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.645 0.070 309.715 ;
    END
  END rd_out_r1[88]
  PIN rd_out_r1[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.065 0.070 310.135 ;
    END
  END rd_out_r1[89]
  PIN rd_out_r1[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.485 0.070 310.555 ;
    END
  END rd_out_r1[90]
  PIN rd_out_r1[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.905 0.070 310.975 ;
    END
  END rd_out_r1[91]
  PIN rd_out_r1[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.325 0.070 311.395 ;
    END
  END rd_out_r1[92]
  PIN rd_out_r1[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.745 0.070 311.815 ;
    END
  END rd_out_r1[93]
  PIN rd_out_r1[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.165 0.070 312.235 ;
    END
  END rd_out_r1[94]
  PIN rd_out_r1[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.585 0.070 312.655 ;
    END
  END rd_out_r1[95]
  PIN rd_out_r1[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.005 0.070 313.075 ;
    END
  END rd_out_r1[96]
  PIN rd_out_r1[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.425 0.070 313.495 ;
    END
  END rd_out_r1[97]
  PIN rd_out_r1[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.845 0.070 313.915 ;
    END
  END rd_out_r1[98]
  PIN rd_out_r1[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.265 0.070 314.335 ;
    END
  END rd_out_r1[99]
  PIN rd_out_r1[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.685 0.070 314.755 ;
    END
  END rd_out_r1[100]
  PIN rd_out_r1[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.105 0.070 315.175 ;
    END
  END rd_out_r1[101]
  PIN rd_out_r1[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.525 0.070 315.595 ;
    END
  END rd_out_r1[102]
  PIN rd_out_r1[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.945 0.070 316.015 ;
    END
  END rd_out_r1[103]
  PIN rd_out_r1[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.365 0.070 316.435 ;
    END
  END rd_out_r1[104]
  PIN rd_out_r1[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.785 0.070 316.855 ;
    END
  END rd_out_r1[105]
  PIN rd_out_r1[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.205 0.070 317.275 ;
    END
  END rd_out_r1[106]
  PIN rd_out_r1[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.625 0.070 317.695 ;
    END
  END rd_out_r1[107]
  PIN rd_out_r1[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.045 0.070 318.115 ;
    END
  END rd_out_r1[108]
  PIN rd_out_r1[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.465 0.070 318.535 ;
    END
  END rd_out_r1[109]
  PIN rd_out_r1[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.885 0.070 318.955 ;
    END
  END rd_out_r1[110]
  PIN rd_out_r1[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 319.305 0.070 319.375 ;
    END
  END rd_out_r1[111]
  PIN rd_out_r1[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 319.725 0.070 319.795 ;
    END
  END rd_out_r1[112]
  PIN rd_out_r1[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.145 0.070 320.215 ;
    END
  END rd_out_r1[113]
  PIN rd_out_r1[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.565 0.070 320.635 ;
    END
  END rd_out_r1[114]
  PIN rd_out_r1[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.985 0.070 321.055 ;
    END
  END rd_out_r1[115]
  PIN rd_out_r1[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.405 0.070 321.475 ;
    END
  END rd_out_r1[116]
  PIN rd_out_r1[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.825 0.070 321.895 ;
    END
  END rd_out_r1[117]
  PIN rd_out_r1[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.245 0.070 322.315 ;
    END
  END rd_out_r1[118]
  PIN rd_out_r1[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.665 0.070 322.735 ;
    END
  END rd_out_r1[119]
  PIN rd_out_r1[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.085 0.070 323.155 ;
    END
  END rd_out_r1[120]
  PIN rd_out_r1[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.505 0.070 323.575 ;
    END
  END rd_out_r1[121]
  PIN rd_out_r1[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.925 0.070 323.995 ;
    END
  END rd_out_r1[122]
  PIN rd_out_r1[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.345 0.070 324.415 ;
    END
  END rd_out_r1[123]
  PIN rd_out_r1[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.765 0.070 324.835 ;
    END
  END rd_out_r1[124]
  PIN rd_out_r1[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.185 0.070 325.255 ;
    END
  END rd_out_r1[125]
  PIN rd_out_r1[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.605 0.070 325.675 ;
    END
  END rd_out_r1[126]
  PIN rd_out_r1[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.025 0.070 326.095 ;
    END
  END rd_out_r1[127]
  PIN rd_out_r1[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.445 0.070 326.515 ;
    END
  END rd_out_r1[128]
  PIN rd_out_r1[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.865 0.070 326.935 ;
    END
  END rd_out_r1[129]
  PIN rd_out_r1[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.285 0.070 327.355 ;
    END
  END rd_out_r1[130]
  PIN rd_out_r1[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.705 0.070 327.775 ;
    END
  END rd_out_r1[131]
  PIN rd_out_r1[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.125 0.070 328.195 ;
    END
  END rd_out_r1[132]
  PIN rd_out_r1[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.545 0.070 328.615 ;
    END
  END rd_out_r1[133]
  PIN rd_out_r1[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.965 0.070 329.035 ;
    END
  END rd_out_r1[134]
  PIN rd_out_r1[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.385 0.070 329.455 ;
    END
  END rd_out_r1[135]
  PIN rd_out_r1[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.805 0.070 329.875 ;
    END
  END rd_out_r1[136]
  PIN rd_out_r1[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 330.225 0.070 330.295 ;
    END
  END rd_out_r1[137]
  PIN rd_out_r1[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 330.645 0.070 330.715 ;
    END
  END rd_out_r1[138]
  PIN rd_out_r1[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.065 0.070 331.135 ;
    END
  END rd_out_r1[139]
  PIN rd_out_r1[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.485 0.070 331.555 ;
    END
  END rd_out_r1[140]
  PIN rd_out_r1[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.905 0.070 331.975 ;
    END
  END rd_out_r1[141]
  PIN rd_out_r1[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.325 0.070 332.395 ;
    END
  END rd_out_r1[142]
  PIN rd_out_r1[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.745 0.070 332.815 ;
    END
  END rd_out_r1[143]
  PIN rd_out_r1[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.165 0.070 333.235 ;
    END
  END rd_out_r1[144]
  PIN rd_out_r1[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.585 0.070 333.655 ;
    END
  END rd_out_r1[145]
  PIN rd_out_r1[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.005 0.070 334.075 ;
    END
  END rd_out_r1[146]
  PIN rd_out_r1[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.425 0.070 334.495 ;
    END
  END rd_out_r1[147]
  PIN rd_out_r1[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.845 0.070 334.915 ;
    END
  END rd_out_r1[148]
  PIN rd_out_r1[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.265 0.070 335.335 ;
    END
  END rd_out_r1[149]
  PIN rd_out_r1[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.685 0.070 335.755 ;
    END
  END rd_out_r1[150]
  PIN rd_out_r1[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.105 0.070 336.175 ;
    END
  END rd_out_r1[151]
  PIN rd_out_r1[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.525 0.070 336.595 ;
    END
  END rd_out_r1[152]
  PIN rd_out_r1[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.945 0.070 337.015 ;
    END
  END rd_out_r1[153]
  PIN rd_out_r1[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.365 0.070 337.435 ;
    END
  END rd_out_r1[154]
  PIN rd_out_r1[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.785 0.070 337.855 ;
    END
  END rd_out_r1[155]
  PIN rd_out_r1[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.205 0.070 338.275 ;
    END
  END rd_out_r1[156]
  PIN rd_out_r1[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.625 0.070 338.695 ;
    END
  END rd_out_r1[157]
  PIN rd_out_r1[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 339.045 0.070 339.115 ;
    END
  END rd_out_r1[158]
  PIN rd_out_r1[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 339.465 0.070 339.535 ;
    END
  END rd_out_r1[159]
  PIN rd_out_r1[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 339.885 0.070 339.955 ;
    END
  END rd_out_r1[160]
  PIN rd_out_r1[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.305 0.070 340.375 ;
    END
  END rd_out_r1[161]
  PIN rd_out_r1[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.725 0.070 340.795 ;
    END
  END rd_out_r1[162]
  PIN rd_out_r1[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.145 0.070 341.215 ;
    END
  END rd_out_r1[163]
  PIN rd_out_r1[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.565 0.070 341.635 ;
    END
  END rd_out_r1[164]
  PIN rd_out_r1[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.985 0.070 342.055 ;
    END
  END rd_out_r1[165]
  PIN rd_out_r1[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.405 0.070 342.475 ;
    END
  END rd_out_r1[166]
  PIN rd_out_r1[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.825 0.070 342.895 ;
    END
  END rd_out_r1[167]
  PIN rd_out_r1[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.245 0.070 343.315 ;
    END
  END rd_out_r1[168]
  PIN rd_out_r1[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.665 0.070 343.735 ;
    END
  END rd_out_r1[169]
  PIN rd_out_r1[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.085 0.070 344.155 ;
    END
  END rd_out_r1[170]
  PIN rd_out_r1[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.505 0.070 344.575 ;
    END
  END rd_out_r1[171]
  PIN rd_out_r1[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.925 0.070 344.995 ;
    END
  END rd_out_r1[172]
  PIN rd_out_r1[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.345 0.070 345.415 ;
    END
  END rd_out_r1[173]
  PIN rd_out_r1[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.765 0.070 345.835 ;
    END
  END rd_out_r1[174]
  PIN rd_out_r1[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.185 0.070 346.255 ;
    END
  END rd_out_r1[175]
  PIN rd_out_r1[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.605 0.070 346.675 ;
    END
  END rd_out_r1[176]
  PIN rd_out_r1[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.025 0.070 347.095 ;
    END
  END rd_out_r1[177]
  PIN rd_out_r1[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.445 0.070 347.515 ;
    END
  END rd_out_r1[178]
  PIN rd_out_r1[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.865 0.070 347.935 ;
    END
  END rd_out_r1[179]
  PIN rd_out_r1[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.285 0.070 348.355 ;
    END
  END rd_out_r1[180]
  PIN rd_out_r1[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.705 0.070 348.775 ;
    END
  END rd_out_r1[181]
  PIN rd_out_r1[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.125 0.070 349.195 ;
    END
  END rd_out_r1[182]
  PIN rd_out_r1[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.545 0.070 349.615 ;
    END
  END rd_out_r1[183]
  PIN rd_out_r1[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.965 0.070 350.035 ;
    END
  END rd_out_r1[184]
  PIN rd_out_r1[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.385 0.070 350.455 ;
    END
  END rd_out_r1[185]
  PIN rd_out_r1[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.805 0.070 350.875 ;
    END
  END rd_out_r1[186]
  PIN rd_out_r1[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.225 0.070 351.295 ;
    END
  END rd_out_r1[187]
  PIN rd_out_r1[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.645 0.070 351.715 ;
    END
  END rd_out_r1[188]
  PIN rd_out_r1[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.065 0.070 352.135 ;
    END
  END rd_out_r1[189]
  PIN rd_out_r1[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.485 0.070 352.555 ;
    END
  END rd_out_r1[190]
  PIN rd_out_r1[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.905 0.070 352.975 ;
    END
  END rd_out_r1[191]
  PIN rd_out_r1[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.325 0.070 353.395 ;
    END
  END rd_out_r1[192]
  PIN rd_out_r1[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.745 0.070 353.815 ;
    END
  END rd_out_r1[193]
  PIN rd_out_r1[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.165 0.070 354.235 ;
    END
  END rd_out_r1[194]
  PIN rd_out_r1[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.585 0.070 354.655 ;
    END
  END rd_out_r1[195]
  PIN rd_out_r1[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.005 0.070 355.075 ;
    END
  END rd_out_r1[196]
  PIN rd_out_r1[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.425 0.070 355.495 ;
    END
  END rd_out_r1[197]
  PIN rd_out_r1[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.845 0.070 355.915 ;
    END
  END rd_out_r1[198]
  PIN rd_out_r1[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.265 0.070 356.335 ;
    END
  END rd_out_r1[199]
  PIN rd_out_r1[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.685 0.070 356.755 ;
    END
  END rd_out_r1[200]
  PIN rd_out_r1[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.105 0.070 357.175 ;
    END
  END rd_out_r1[201]
  PIN rd_out_r1[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.525 0.070 357.595 ;
    END
  END rd_out_r1[202]
  PIN rd_out_r1[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.945 0.070 358.015 ;
    END
  END rd_out_r1[203]
  PIN rd_out_r1[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.365 0.070 358.435 ;
    END
  END rd_out_r1[204]
  PIN rd_out_r1[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.785 0.070 358.855 ;
    END
  END rd_out_r1[205]
  PIN rd_out_r1[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.205 0.070 359.275 ;
    END
  END rd_out_r1[206]
  PIN rd_out_r1[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.625 0.070 359.695 ;
    END
  END rd_out_r1[207]
  PIN rd_out_r1[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.045 0.070 360.115 ;
    END
  END rd_out_r1[208]
  PIN rd_out_r1[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.465 0.070 360.535 ;
    END
  END rd_out_r1[209]
  PIN rd_out_r1[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.885 0.070 360.955 ;
    END
  END rd_out_r1[210]
  PIN rd_out_r1[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 361.305 0.070 361.375 ;
    END
  END rd_out_r1[211]
  PIN rd_out_r1[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 361.725 0.070 361.795 ;
    END
  END rd_out_r1[212]
  PIN rd_out_r1[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.145 0.070 362.215 ;
    END
  END rd_out_r1[213]
  PIN rd_out_r1[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.565 0.070 362.635 ;
    END
  END rd_out_r1[214]
  PIN rd_out_r1[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.985 0.070 363.055 ;
    END
  END rd_out_r1[215]
  PIN rd_out_r1[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.405 0.070 363.475 ;
    END
  END rd_out_r1[216]
  PIN rd_out_r1[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.825 0.070 363.895 ;
    END
  END rd_out_r1[217]
  PIN rd_out_r1[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.245 0.070 364.315 ;
    END
  END rd_out_r1[218]
  PIN rd_out_r1[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.665 0.070 364.735 ;
    END
  END rd_out_r1[219]
  PIN rd_out_r1[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.085 0.070 365.155 ;
    END
  END rd_out_r1[220]
  PIN rd_out_r1[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.505 0.070 365.575 ;
    END
  END rd_out_r1[221]
  PIN rd_out_r1[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.925 0.070 365.995 ;
    END
  END rd_out_r1[222]
  PIN rd_out_r1[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 366.345 0.070 366.415 ;
    END
  END rd_out_r1[223]
  PIN rd_out_r1[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 366.765 0.070 366.835 ;
    END
  END rd_out_r1[224]
  PIN rd_out_r1[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.185 0.070 367.255 ;
    END
  END rd_out_r1[225]
  PIN rd_out_r1[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.605 0.070 367.675 ;
    END
  END rd_out_r1[226]
  PIN rd_out_r1[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.025 0.070 368.095 ;
    END
  END rd_out_r1[227]
  PIN rd_out_r1[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.445 0.070 368.515 ;
    END
  END rd_out_r1[228]
  PIN rd_out_r1[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.865 0.070 368.935 ;
    END
  END rd_out_r1[229]
  PIN rd_out_r1[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.285 0.070 369.355 ;
    END
  END rd_out_r1[230]
  PIN rd_out_r1[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.705 0.070 369.775 ;
    END
  END rd_out_r1[231]
  PIN rd_out_r1[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.125 0.070 370.195 ;
    END
  END rd_out_r1[232]
  PIN rd_out_r1[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.545 0.070 370.615 ;
    END
  END rd_out_r1[233]
  PIN rd_out_r1[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.965 0.070 371.035 ;
    END
  END rd_out_r1[234]
  PIN rd_out_r1[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 371.385 0.070 371.455 ;
    END
  END rd_out_r1[235]
  PIN rd_out_r1[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 371.805 0.070 371.875 ;
    END
  END rd_out_r1[236]
  PIN rd_out_r1[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.225 0.070 372.295 ;
    END
  END rd_out_r1[237]
  PIN rd_out_r1[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.645 0.070 372.715 ;
    END
  END rd_out_r1[238]
  PIN rd_out_r1[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.065 0.070 373.135 ;
    END
  END rd_out_r1[239]
  PIN rd_out_r1[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.485 0.070 373.555 ;
    END
  END rd_out_r1[240]
  PIN rd_out_r1[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.905 0.070 373.975 ;
    END
  END rd_out_r1[241]
  PIN rd_out_r1[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.325 0.070 374.395 ;
    END
  END rd_out_r1[242]
  PIN rd_out_r1[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.745 0.070 374.815 ;
    END
  END rd_out_r1[243]
  PIN rd_out_r1[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 375.165 0.070 375.235 ;
    END
  END rd_out_r1[244]
  PIN rd_out_r1[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 375.585 0.070 375.655 ;
    END
  END rd_out_r1[245]
  PIN rd_out_r1[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.005 0.070 376.075 ;
    END
  END rd_out_r1[246]
  PIN rd_out_r1[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.425 0.070 376.495 ;
    END
  END rd_out_r1[247]
  PIN rd_out_r1[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.845 0.070 376.915 ;
    END
  END rd_out_r1[248]
  PIN rd_out_r1[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.265 0.070 377.335 ;
    END
  END rd_out_r1[249]
  PIN rd_out_r1[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.685 0.070 377.755 ;
    END
  END rd_out_r1[250]
  PIN rd_out_r1[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.105 0.070 378.175 ;
    END
  END rd_out_r1[251]
  PIN rd_out_r1[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.525 0.070 378.595 ;
    END
  END rd_out_r1[252]
  PIN rd_out_r1[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.945 0.070 379.015 ;
    END
  END rd_out_r1[253]
  PIN rd_out_r1[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.365 0.070 379.435 ;
    END
  END rd_out_r1[254]
  PIN rd_out_r1[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.785 0.070 379.855 ;
    END
  END rd_out_r1[255]
  PIN rd_out_r1[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 380.205 0.070 380.275 ;
    END
  END rd_out_r1[256]
  PIN rd_out_r1[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 380.625 0.070 380.695 ;
    END
  END rd_out_r1[257]
  PIN rd_out_r1[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.045 0.070 381.115 ;
    END
  END rd_out_r1[258]
  PIN rd_out_r1[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.465 0.070 381.535 ;
    END
  END rd_out_r1[259]
  PIN rd_out_r1[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.885 0.070 381.955 ;
    END
  END rd_out_r1[260]
  PIN rd_out_r1[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 382.305 0.070 382.375 ;
    END
  END rd_out_r1[261]
  PIN rd_out_r1[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 382.725 0.070 382.795 ;
    END
  END rd_out_r1[262]
  PIN rd_out_r1[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.145 0.070 383.215 ;
    END
  END rd_out_r1[263]
  PIN rd_out_r1[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.565 0.070 383.635 ;
    END
  END rd_out_r1[264]
  PIN rd_out_r1[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.985 0.070 384.055 ;
    END
  END rd_out_r1[265]
  PIN rd_out_r1[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.405 0.070 384.475 ;
    END
  END rd_out_r1[266]
  PIN rd_out_r1[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.825 0.070 384.895 ;
    END
  END rd_out_r1[267]
  PIN rd_out_r1[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.245 0.070 385.315 ;
    END
  END rd_out_r1[268]
  PIN rd_out_r1[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.665 0.070 385.735 ;
    END
  END rd_out_r1[269]
  PIN rd_out_r1[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.085 0.070 386.155 ;
    END
  END rd_out_r1[270]
  PIN rd_out_r1[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.505 0.070 386.575 ;
    END
  END rd_out_r1[271]
  PIN rd_out_r1[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.925 0.070 386.995 ;
    END
  END rd_out_r1[272]
  PIN rd_out_r1[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.345 0.070 387.415 ;
    END
  END rd_out_r1[273]
  PIN rd_out_r1[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.765 0.070 387.835 ;
    END
  END rd_out_r1[274]
  PIN rd_out_r1[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.185 0.070 388.255 ;
    END
  END rd_out_r1[275]
  PIN rd_out_r1[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.605 0.070 388.675 ;
    END
  END rd_out_r1[276]
  PIN rd_out_r1[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 389.025 0.070 389.095 ;
    END
  END rd_out_r1[277]
  PIN rd_out_r1[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 389.445 0.070 389.515 ;
    END
  END rd_out_r1[278]
  PIN rd_out_r1[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 389.865 0.070 389.935 ;
    END
  END rd_out_r1[279]
  PIN rd_out_r1[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.285 0.070 390.355 ;
    END
  END rd_out_r1[280]
  PIN rd_out_r1[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.705 0.070 390.775 ;
    END
  END rd_out_r1[281]
  PIN rd_out_r1[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.125 0.070 391.195 ;
    END
  END rd_out_r1[282]
  PIN rd_out_r1[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.545 0.070 391.615 ;
    END
  END rd_out_r1[283]
  PIN rd_out_r1[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.965 0.070 392.035 ;
    END
  END rd_out_r1[284]
  PIN rd_out_r1[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.385 0.070 392.455 ;
    END
  END rd_out_r1[285]
  PIN rd_out_r1[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.805 0.070 392.875 ;
    END
  END rd_out_r1[286]
  PIN rd_out_r1[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.225 0.070 393.295 ;
    END
  END rd_out_r1[287]
  PIN rd_out_r1[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.645 0.070 393.715 ;
    END
  END rd_out_r1[288]
  PIN rd_out_r1[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.065 0.070 394.135 ;
    END
  END rd_out_r1[289]
  PIN rd_out_r1[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.485 0.070 394.555 ;
    END
  END rd_out_r1[290]
  PIN rd_out_r1[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.905 0.070 394.975 ;
    END
  END rd_out_r1[291]
  PIN rd_out_r1[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.325 0.070 395.395 ;
    END
  END rd_out_r1[292]
  PIN rd_out_r1[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.745 0.070 395.815 ;
    END
  END rd_out_r1[293]
  PIN rd_out_r1[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.165 0.070 396.235 ;
    END
  END rd_out_r1[294]
  PIN rd_out_r1[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.585 0.070 396.655 ;
    END
  END rd_out_r1[295]
  PIN rd_out_r1[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.005 0.070 397.075 ;
    END
  END rd_out_r1[296]
  PIN rd_out_r1[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.425 0.070 397.495 ;
    END
  END rd_out_r1[297]
  PIN rd_out_r1[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.845 0.070 397.915 ;
    END
  END rd_out_r1[298]
  PIN rd_out_r1[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.265 0.070 398.335 ;
    END
  END rd_out_r1[299]
  PIN rd_out_r1[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.685 0.070 398.755 ;
    END
  END rd_out_r1[300]
  PIN rd_out_r1[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.105 0.070 399.175 ;
    END
  END rd_out_r1[301]
  PIN rd_out_r1[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.525 0.070 399.595 ;
    END
  END rd_out_r1[302]
  PIN rd_out_r1[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.945 0.070 400.015 ;
    END
  END rd_out_r1[303]
  PIN rd_out_r1[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 400.365 0.070 400.435 ;
    END
  END rd_out_r1[304]
  PIN rd_out_r1[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 400.785 0.070 400.855 ;
    END
  END rd_out_r1[305]
  PIN rd_out_r1[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 401.205 0.070 401.275 ;
    END
  END rd_out_r1[306]
  PIN rd_out_r1[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 401.625 0.070 401.695 ;
    END
  END rd_out_r1[307]
  PIN rd_out_r1[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 402.045 0.070 402.115 ;
    END
  END rd_out_r1[308]
  PIN rd_out_r1[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 402.465 0.070 402.535 ;
    END
  END rd_out_r1[309]
  PIN rd_out_r1[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 402.885 0.070 402.955 ;
    END
  END rd_out_r1[310]
  PIN rd_out_r1[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 403.305 0.070 403.375 ;
    END
  END rd_out_r1[311]
  PIN rd_out_r1[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 403.725 0.070 403.795 ;
    END
  END rd_out_r1[312]
  PIN rd_out_r1[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 404.145 0.070 404.215 ;
    END
  END rd_out_r1[313]
  PIN rd_out_r1[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 404.565 0.070 404.635 ;
    END
  END rd_out_r1[314]
  PIN rd_out_r1[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 404.985 0.070 405.055 ;
    END
  END rd_out_r1[315]
  PIN rd_out_r1[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 405.405 0.070 405.475 ;
    END
  END rd_out_r1[316]
  PIN rd_out_r1[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 405.825 0.070 405.895 ;
    END
  END rd_out_r1[317]
  PIN rd_out_r1[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 406.245 0.070 406.315 ;
    END
  END rd_out_r1[318]
  PIN rd_out_r1[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 406.665 0.070 406.735 ;
    END
  END rd_out_r1[319]
  PIN rd_out_r1[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 407.085 0.070 407.155 ;
    END
  END rd_out_r1[320]
  PIN rd_out_r1[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 407.505 0.070 407.575 ;
    END
  END rd_out_r1[321]
  PIN rd_out_r1[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 407.925 0.070 407.995 ;
    END
  END rd_out_r1[322]
  PIN rd_out_r1[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 408.345 0.070 408.415 ;
    END
  END rd_out_r1[323]
  PIN rd_out_r1[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 408.765 0.070 408.835 ;
    END
  END rd_out_r1[324]
  PIN rd_out_r1[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 409.185 0.070 409.255 ;
    END
  END rd_out_r1[325]
  PIN rd_out_r1[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 409.605 0.070 409.675 ;
    END
  END rd_out_r1[326]
  PIN rd_out_r1[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 410.025 0.070 410.095 ;
    END
  END rd_out_r1[327]
  PIN rd_out_r1[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 410.445 0.070 410.515 ;
    END
  END rd_out_r1[328]
  PIN rd_out_r1[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 410.865 0.070 410.935 ;
    END
  END rd_out_r1[329]
  PIN rd_out_r1[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 411.285 0.070 411.355 ;
    END
  END rd_out_r1[330]
  PIN rd_out_r1[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 411.705 0.070 411.775 ;
    END
  END rd_out_r1[331]
  PIN rd_out_r1[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 412.125 0.070 412.195 ;
    END
  END rd_out_r1[332]
  PIN rd_out_r1[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 412.545 0.070 412.615 ;
    END
  END rd_out_r1[333]
  PIN rd_out_r1[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 412.965 0.070 413.035 ;
    END
  END rd_out_r1[334]
  PIN rd_out_r1[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 413.385 0.070 413.455 ;
    END
  END rd_out_r1[335]
  PIN rd_out_r1[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 413.805 0.070 413.875 ;
    END
  END rd_out_r1[336]
  PIN rd_out_r1[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 414.225 0.070 414.295 ;
    END
  END rd_out_r1[337]
  PIN rd_out_r1[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 414.645 0.070 414.715 ;
    END
  END rd_out_r1[338]
  PIN rd_out_r1[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 415.065 0.070 415.135 ;
    END
  END rd_out_r1[339]
  PIN rd_out_r1[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 415.485 0.070 415.555 ;
    END
  END rd_out_r1[340]
  PIN rd_out_r1[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 415.905 0.070 415.975 ;
    END
  END rd_out_r1[341]
  PIN rd_out_r1[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 416.325 0.070 416.395 ;
    END
  END rd_out_r1[342]
  PIN rd_out_r1[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 416.745 0.070 416.815 ;
    END
  END rd_out_r1[343]
  PIN rd_out_r1[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 417.165 0.070 417.235 ;
    END
  END rd_out_r1[344]
  PIN rd_out_r1[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 417.585 0.070 417.655 ;
    END
  END rd_out_r1[345]
  PIN rd_out_r1[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 418.005 0.070 418.075 ;
    END
  END rd_out_r1[346]
  PIN rd_out_r1[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 418.425 0.070 418.495 ;
    END
  END rd_out_r1[347]
  PIN rd_out_r1[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 418.845 0.070 418.915 ;
    END
  END rd_out_r1[348]
  PIN rd_out_r1[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 419.265 0.070 419.335 ;
    END
  END rd_out_r1[349]
  PIN rd_out_r1[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 419.685 0.070 419.755 ;
    END
  END rd_out_r1[350]
  PIN rd_out_r1[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 420.105 0.070 420.175 ;
    END
  END rd_out_r1[351]
  PIN rd_out_r1[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 420.525 0.070 420.595 ;
    END
  END rd_out_r1[352]
  PIN rd_out_r1[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 420.945 0.070 421.015 ;
    END
  END rd_out_r1[353]
  PIN rd_out_r1[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 421.365 0.070 421.435 ;
    END
  END rd_out_r1[354]
  PIN rd_out_r1[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 421.785 0.070 421.855 ;
    END
  END rd_out_r1[355]
  PIN rd_out_r1[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 422.205 0.070 422.275 ;
    END
  END rd_out_r1[356]
  PIN rd_out_r1[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 422.625 0.070 422.695 ;
    END
  END rd_out_r1[357]
  PIN rd_out_r1[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 423.045 0.070 423.115 ;
    END
  END rd_out_r1[358]
  PIN rd_out_r1[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 423.465 0.070 423.535 ;
    END
  END rd_out_r1[359]
  PIN rd_out_r1[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 423.885 0.070 423.955 ;
    END
  END rd_out_r1[360]
  PIN rd_out_r1[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 424.305 0.070 424.375 ;
    END
  END rd_out_r1[361]
  PIN rd_out_r1[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 424.725 0.070 424.795 ;
    END
  END rd_out_r1[362]
  PIN rd_out_r1[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 425.145 0.070 425.215 ;
    END
  END rd_out_r1[363]
  PIN rd_out_r1[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 425.565 0.070 425.635 ;
    END
  END rd_out_r1[364]
  PIN rd_out_r1[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 425.985 0.070 426.055 ;
    END
  END rd_out_r1[365]
  PIN rd_out_r1[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 426.405 0.070 426.475 ;
    END
  END rd_out_r1[366]
  PIN rd_out_r1[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 426.825 0.070 426.895 ;
    END
  END rd_out_r1[367]
  PIN rd_out_r1[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 427.245 0.070 427.315 ;
    END
  END rd_out_r1[368]
  PIN rd_out_r1[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 427.665 0.070 427.735 ;
    END
  END rd_out_r1[369]
  PIN rd_out_r1[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 428.085 0.070 428.155 ;
    END
  END rd_out_r1[370]
  PIN rd_out_r1[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 428.505 0.070 428.575 ;
    END
  END rd_out_r1[371]
  PIN rd_out_r1[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 428.925 0.070 428.995 ;
    END
  END rd_out_r1[372]
  PIN rd_out_r1[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 429.345 0.070 429.415 ;
    END
  END rd_out_r1[373]
  PIN rd_out_r1[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 429.765 0.070 429.835 ;
    END
  END rd_out_r1[374]
  PIN rd_out_r1[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 430.185 0.070 430.255 ;
    END
  END rd_out_r1[375]
  PIN rd_out_r1[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 430.605 0.070 430.675 ;
    END
  END rd_out_r1[376]
  PIN rd_out_r1[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 431.025 0.070 431.095 ;
    END
  END rd_out_r1[377]
  PIN rd_out_r1[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 431.445 0.070 431.515 ;
    END
  END rd_out_r1[378]
  PIN rd_out_r1[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 431.865 0.070 431.935 ;
    END
  END rd_out_r1[379]
  PIN rd_out_r1[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 432.285 0.070 432.355 ;
    END
  END rd_out_r1[380]
  PIN rd_out_r1[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 432.705 0.070 432.775 ;
    END
  END rd_out_r1[381]
  PIN rd_out_r1[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 433.125 0.070 433.195 ;
    END
  END rd_out_r1[382]
  PIN rd_out_r1[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 433.545 0.070 433.615 ;
    END
  END rd_out_r1[383]
  PIN rd_out_r1[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 433.965 0.070 434.035 ;
    END
  END rd_out_r1[384]
  PIN rd_out_r1[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 434.385 0.070 434.455 ;
    END
  END rd_out_r1[385]
  PIN rd_out_r1[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 434.805 0.070 434.875 ;
    END
  END rd_out_r1[386]
  PIN rd_out_r1[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 435.225 0.070 435.295 ;
    END
  END rd_out_r1[387]
  PIN rd_out_r1[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 435.645 0.070 435.715 ;
    END
  END rd_out_r1[388]
  PIN rd_out_r1[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 436.065 0.070 436.135 ;
    END
  END rd_out_r1[389]
  PIN rd_out_r1[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 436.485 0.070 436.555 ;
    END
  END rd_out_r1[390]
  PIN rd_out_r1[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 436.905 0.070 436.975 ;
    END
  END rd_out_r1[391]
  PIN rd_out_r1[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 437.325 0.070 437.395 ;
    END
  END rd_out_r1[392]
  PIN rd_out_r1[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 437.745 0.070 437.815 ;
    END
  END rd_out_r1[393]
  PIN rd_out_r1[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 438.165 0.070 438.235 ;
    END
  END rd_out_r1[394]
  PIN rd_out_r1[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 438.585 0.070 438.655 ;
    END
  END rd_out_r1[395]
  PIN rd_out_r1[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 439.005 0.070 439.075 ;
    END
  END rd_out_r1[396]
  PIN rd_out_r1[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 439.425 0.070 439.495 ;
    END
  END rd_out_r1[397]
  PIN rd_out_r1[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 439.845 0.070 439.915 ;
    END
  END rd_out_r1[398]
  PIN rd_out_r1[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 440.265 0.070 440.335 ;
    END
  END rd_out_r1[399]
  PIN rd_out_r1[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 440.685 0.070 440.755 ;
    END
  END rd_out_r1[400]
  PIN rd_out_r1[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 441.105 0.070 441.175 ;
    END
  END rd_out_r1[401]
  PIN rd_out_r1[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 441.525 0.070 441.595 ;
    END
  END rd_out_r1[402]
  PIN rd_out_r1[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 441.945 0.070 442.015 ;
    END
  END rd_out_r1[403]
  PIN rd_out_r1[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 442.365 0.070 442.435 ;
    END
  END rd_out_r1[404]
  PIN rd_out_r1[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 442.785 0.070 442.855 ;
    END
  END rd_out_r1[405]
  PIN rd_out_r1[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 443.205 0.070 443.275 ;
    END
  END rd_out_r1[406]
  PIN rd_out_r1[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 443.625 0.070 443.695 ;
    END
  END rd_out_r1[407]
  PIN rd_out_r1[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 444.045 0.070 444.115 ;
    END
  END rd_out_r1[408]
  PIN rd_out_r1[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 444.465 0.070 444.535 ;
    END
  END rd_out_r1[409]
  PIN rd_out_r1[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 444.885 0.070 444.955 ;
    END
  END rd_out_r1[410]
  PIN rd_out_r1[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 445.305 0.070 445.375 ;
    END
  END rd_out_r1[411]
  PIN rd_out_r1[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 445.725 0.070 445.795 ;
    END
  END rd_out_r1[412]
  PIN rd_out_r1[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 446.145 0.070 446.215 ;
    END
  END rd_out_r1[413]
  PIN rd_out_r1[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 446.565 0.070 446.635 ;
    END
  END rd_out_r1[414]
  PIN rd_out_r1[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 446.985 0.070 447.055 ;
    END
  END rd_out_r1[415]
  PIN rd_out_r1[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 447.405 0.070 447.475 ;
    END
  END rd_out_r1[416]
  PIN rd_out_r1[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 447.825 0.070 447.895 ;
    END
  END rd_out_r1[417]
  PIN rd_out_r1[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 448.245 0.070 448.315 ;
    END
  END rd_out_r1[418]
  PIN rd_out_r1[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 448.665 0.070 448.735 ;
    END
  END rd_out_r1[419]
  PIN rd_out_r1[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 449.085 0.070 449.155 ;
    END
  END rd_out_r1[420]
  PIN rd_out_r1[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 449.505 0.070 449.575 ;
    END
  END rd_out_r1[421]
  PIN rd_out_r1[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 449.925 0.070 449.995 ;
    END
  END rd_out_r1[422]
  PIN rd_out_r1[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 450.345 0.070 450.415 ;
    END
  END rd_out_r1[423]
  PIN rd_out_r1[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 450.765 0.070 450.835 ;
    END
  END rd_out_r1[424]
  PIN rd_out_r1[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 451.185 0.070 451.255 ;
    END
  END rd_out_r1[425]
  PIN rd_out_r1[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 451.605 0.070 451.675 ;
    END
  END rd_out_r1[426]
  PIN rd_out_r1[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 452.025 0.070 452.095 ;
    END
  END rd_out_r1[427]
  PIN rd_out_r1[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 452.445 0.070 452.515 ;
    END
  END rd_out_r1[428]
  PIN rd_out_r1[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 452.865 0.070 452.935 ;
    END
  END rd_out_r1[429]
  PIN rd_out_r1[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 453.285 0.070 453.355 ;
    END
  END rd_out_r1[430]
  PIN rd_out_r1[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 453.705 0.070 453.775 ;
    END
  END rd_out_r1[431]
  PIN rd_out_r1[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 454.125 0.070 454.195 ;
    END
  END rd_out_r1[432]
  PIN rd_out_r1[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 454.545 0.070 454.615 ;
    END
  END rd_out_r1[433]
  PIN rd_out_r1[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 454.965 0.070 455.035 ;
    END
  END rd_out_r1[434]
  PIN rd_out_r1[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 455.385 0.070 455.455 ;
    END
  END rd_out_r1[435]
  PIN rd_out_r1[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 455.805 0.070 455.875 ;
    END
  END rd_out_r1[436]
  PIN rd_out_r1[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 456.225 0.070 456.295 ;
    END
  END rd_out_r1[437]
  PIN rd_out_r1[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 456.645 0.070 456.715 ;
    END
  END rd_out_r1[438]
  PIN rd_out_r1[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 457.065 0.070 457.135 ;
    END
  END rd_out_r1[439]
  PIN rd_out_r1[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 457.485 0.070 457.555 ;
    END
  END rd_out_r1[440]
  PIN rd_out_r1[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 457.905 0.070 457.975 ;
    END
  END rd_out_r1[441]
  PIN rd_out_r1[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 458.325 0.070 458.395 ;
    END
  END rd_out_r1[442]
  PIN rd_out_r1[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 458.745 0.070 458.815 ;
    END
  END rd_out_r1[443]
  PIN rd_out_r1[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 459.165 0.070 459.235 ;
    END
  END rd_out_r1[444]
  PIN rd_out_r1[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 459.585 0.070 459.655 ;
    END
  END rd_out_r1[445]
  PIN rd_out_r1[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 460.005 0.070 460.075 ;
    END
  END rd_out_r1[446]
  PIN rd_out_r1[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 460.425 0.070 460.495 ;
    END
  END rd_out_r1[447]
  PIN rd_out_r1[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 460.845 0.070 460.915 ;
    END
  END rd_out_r1[448]
  PIN rd_out_r1[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 461.265 0.070 461.335 ;
    END
  END rd_out_r1[449]
  PIN rd_out_r1[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 461.685 0.070 461.755 ;
    END
  END rd_out_r1[450]
  PIN rd_out_r1[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 462.105 0.070 462.175 ;
    END
  END rd_out_r1[451]
  PIN rd_out_r1[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 462.525 0.070 462.595 ;
    END
  END rd_out_r1[452]
  PIN rd_out_r1[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 462.945 0.070 463.015 ;
    END
  END rd_out_r1[453]
  PIN rd_out_r1[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 463.365 0.070 463.435 ;
    END
  END rd_out_r1[454]
  PIN rd_out_r1[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 463.785 0.070 463.855 ;
    END
  END rd_out_r1[455]
  PIN rd_out_r1[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 464.205 0.070 464.275 ;
    END
  END rd_out_r1[456]
  PIN rd_out_r1[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 464.625 0.070 464.695 ;
    END
  END rd_out_r1[457]
  PIN rd_out_r1[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 465.045 0.070 465.115 ;
    END
  END rd_out_r1[458]
  PIN rd_out_r1[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 465.465 0.070 465.535 ;
    END
  END rd_out_r1[459]
  PIN rd_out_r1[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 465.885 0.070 465.955 ;
    END
  END rd_out_r1[460]
  PIN rd_out_r1[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 466.305 0.070 466.375 ;
    END
  END rd_out_r1[461]
  PIN rd_out_r1[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 466.725 0.070 466.795 ;
    END
  END rd_out_r1[462]
  PIN rd_out_r1[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 467.145 0.070 467.215 ;
    END
  END rd_out_r1[463]
  PIN rd_out_r1[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 467.565 0.070 467.635 ;
    END
  END rd_out_r1[464]
  PIN rd_out_r1[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 467.985 0.070 468.055 ;
    END
  END rd_out_r1[465]
  PIN rd_out_r1[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 468.405 0.070 468.475 ;
    END
  END rd_out_r1[466]
  PIN rd_out_r1[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 468.825 0.070 468.895 ;
    END
  END rd_out_r1[467]
  PIN rd_out_r1[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 469.245 0.070 469.315 ;
    END
  END rd_out_r1[468]
  PIN rd_out_r1[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 469.665 0.070 469.735 ;
    END
  END rd_out_r1[469]
  PIN rd_out_r1[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 470.085 0.070 470.155 ;
    END
  END rd_out_r1[470]
  PIN rd_out_r1[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 470.505 0.070 470.575 ;
    END
  END rd_out_r1[471]
  PIN rd_out_r1[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 470.925 0.070 470.995 ;
    END
  END rd_out_r1[472]
  PIN rd_out_r1[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 471.345 0.070 471.415 ;
    END
  END rd_out_r1[473]
  PIN rd_out_r1[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 471.765 0.070 471.835 ;
    END
  END rd_out_r1[474]
  PIN rd_out_r1[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 472.185 0.070 472.255 ;
    END
  END rd_out_r1[475]
  PIN rd_out_r1[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 472.605 0.070 472.675 ;
    END
  END rd_out_r1[476]
  PIN rd_out_r1[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 473.025 0.070 473.095 ;
    END
  END rd_out_r1[477]
  PIN rd_out_r1[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 473.445 0.070 473.515 ;
    END
  END rd_out_r1[478]
  PIN rd_out_r1[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 473.865 0.070 473.935 ;
    END
  END rd_out_r1[479]
  PIN rd_out_r1[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 474.285 0.070 474.355 ;
    END
  END rd_out_r1[480]
  PIN rd_out_r1[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 474.705 0.070 474.775 ;
    END
  END rd_out_r1[481]
  PIN rd_out_r1[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 475.125 0.070 475.195 ;
    END
  END rd_out_r1[482]
  PIN rd_out_r1[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 475.545 0.070 475.615 ;
    END
  END rd_out_r1[483]
  PIN rd_out_r1[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 475.965 0.070 476.035 ;
    END
  END rd_out_r1[484]
  PIN rd_out_r1[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 476.385 0.070 476.455 ;
    END
  END rd_out_r1[485]
  PIN rd_out_r1[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 476.805 0.070 476.875 ;
    END
  END rd_out_r1[486]
  PIN rd_out_r1[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 477.225 0.070 477.295 ;
    END
  END rd_out_r1[487]
  PIN rd_out_r1[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 477.645 0.070 477.715 ;
    END
  END rd_out_r1[488]
  PIN rd_out_r1[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 478.065 0.070 478.135 ;
    END
  END rd_out_r1[489]
  PIN rd_out_r1[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 478.485 0.070 478.555 ;
    END
  END rd_out_r1[490]
  PIN rd_out_r1[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 478.905 0.070 478.975 ;
    END
  END rd_out_r1[491]
  PIN rd_out_r1[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 479.325 0.070 479.395 ;
    END
  END rd_out_r1[492]
  PIN rd_out_r1[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 479.745 0.070 479.815 ;
    END
  END rd_out_r1[493]
  PIN rd_out_r1[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 480.165 0.070 480.235 ;
    END
  END rd_out_r1[494]
  PIN rd_out_r1[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 480.585 0.070 480.655 ;
    END
  END rd_out_r1[495]
  PIN rd_out_r1[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 481.005 0.070 481.075 ;
    END
  END rd_out_r1[496]
  PIN rd_out_r1[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 481.425 0.070 481.495 ;
    END
  END rd_out_r1[497]
  PIN rd_out_r1[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 481.845 0.070 481.915 ;
    END
  END rd_out_r1[498]
  PIN rd_out_r1[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 482.265 0.070 482.335 ;
    END
  END rd_out_r1[499]
  PIN rd_out_r1[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 482.685 0.070 482.755 ;
    END
  END rd_out_r1[500]
  PIN rd_out_r1[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 483.105 0.070 483.175 ;
    END
  END rd_out_r1[501]
  PIN rd_out_r1[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 483.525 0.070 483.595 ;
    END
  END rd_out_r1[502]
  PIN rd_out_r1[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 483.945 0.070 484.015 ;
    END
  END rd_out_r1[503]
  PIN rd_out_r1[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 484.365 0.070 484.435 ;
    END
  END rd_out_r1[504]
  PIN rd_out_r1[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 484.785 0.070 484.855 ;
    END
  END rd_out_r1[505]
  PIN rd_out_r1[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 485.205 0.070 485.275 ;
    END
  END rd_out_r1[506]
  PIN rd_out_r1[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 485.625 0.070 485.695 ;
    END
  END rd_out_r1[507]
  PIN rd_out_r1[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 486.045 0.070 486.115 ;
    END
  END rd_out_r1[508]
  PIN rd_out_r1[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 486.465 0.070 486.535 ;
    END
  END rd_out_r1[509]
  PIN rd_out_r1[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 486.885 0.070 486.955 ;
    END
  END rd_out_r1[510]
  PIN rd_out_r1[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 487.305 0.070 487.375 ;
    END
  END rd_out_r1[511]
  PIN wd_in_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 515.865 0.070 515.935 ;
    END
  END wd_in_w1[0]
  PIN wd_in_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.285 0.070 516.355 ;
    END
  END wd_in_w1[1]
  PIN wd_in_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.705 0.070 516.775 ;
    END
  END wd_in_w1[2]
  PIN wd_in_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.125 0.070 517.195 ;
    END
  END wd_in_w1[3]
  PIN wd_in_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.545 0.070 517.615 ;
    END
  END wd_in_w1[4]
  PIN wd_in_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.965 0.070 518.035 ;
    END
  END wd_in_w1[5]
  PIN wd_in_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.385 0.070 518.455 ;
    END
  END wd_in_w1[6]
  PIN wd_in_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.805 0.070 518.875 ;
    END
  END wd_in_w1[7]
  PIN wd_in_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.225 0.070 519.295 ;
    END
  END wd_in_w1[8]
  PIN wd_in_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.645 0.070 519.715 ;
    END
  END wd_in_w1[9]
  PIN wd_in_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.065 0.070 520.135 ;
    END
  END wd_in_w1[10]
  PIN wd_in_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.485 0.070 520.555 ;
    END
  END wd_in_w1[11]
  PIN wd_in_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.905 0.070 520.975 ;
    END
  END wd_in_w1[12]
  PIN wd_in_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.325 0.070 521.395 ;
    END
  END wd_in_w1[13]
  PIN wd_in_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.745 0.070 521.815 ;
    END
  END wd_in_w1[14]
  PIN wd_in_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.165 0.070 522.235 ;
    END
  END wd_in_w1[15]
  PIN wd_in_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.585 0.070 522.655 ;
    END
  END wd_in_w1[16]
  PIN wd_in_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.005 0.070 523.075 ;
    END
  END wd_in_w1[17]
  PIN wd_in_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.425 0.070 523.495 ;
    END
  END wd_in_w1[18]
  PIN wd_in_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.845 0.070 523.915 ;
    END
  END wd_in_w1[19]
  PIN wd_in_w1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.265 0.070 524.335 ;
    END
  END wd_in_w1[20]
  PIN wd_in_w1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.685 0.070 524.755 ;
    END
  END wd_in_w1[21]
  PIN wd_in_w1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.105 0.070 525.175 ;
    END
  END wd_in_w1[22]
  PIN wd_in_w1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.525 0.070 525.595 ;
    END
  END wd_in_w1[23]
  PIN wd_in_w1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.945 0.070 526.015 ;
    END
  END wd_in_w1[24]
  PIN wd_in_w1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.365 0.070 526.435 ;
    END
  END wd_in_w1[25]
  PIN wd_in_w1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.785 0.070 526.855 ;
    END
  END wd_in_w1[26]
  PIN wd_in_w1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.205 0.070 527.275 ;
    END
  END wd_in_w1[27]
  PIN wd_in_w1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.625 0.070 527.695 ;
    END
  END wd_in_w1[28]
  PIN wd_in_w1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.045 0.070 528.115 ;
    END
  END wd_in_w1[29]
  PIN wd_in_w1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.465 0.070 528.535 ;
    END
  END wd_in_w1[30]
  PIN wd_in_w1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.885 0.070 528.955 ;
    END
  END wd_in_w1[31]
  PIN wd_in_w1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.305 0.070 529.375 ;
    END
  END wd_in_w1[32]
  PIN wd_in_w1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.725 0.070 529.795 ;
    END
  END wd_in_w1[33]
  PIN wd_in_w1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.145 0.070 530.215 ;
    END
  END wd_in_w1[34]
  PIN wd_in_w1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.565 0.070 530.635 ;
    END
  END wd_in_w1[35]
  PIN wd_in_w1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.985 0.070 531.055 ;
    END
  END wd_in_w1[36]
  PIN wd_in_w1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.405 0.070 531.475 ;
    END
  END wd_in_w1[37]
  PIN wd_in_w1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.825 0.070 531.895 ;
    END
  END wd_in_w1[38]
  PIN wd_in_w1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.245 0.070 532.315 ;
    END
  END wd_in_w1[39]
  PIN wd_in_w1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.665 0.070 532.735 ;
    END
  END wd_in_w1[40]
  PIN wd_in_w1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.085 0.070 533.155 ;
    END
  END wd_in_w1[41]
  PIN wd_in_w1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.505 0.070 533.575 ;
    END
  END wd_in_w1[42]
  PIN wd_in_w1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.925 0.070 533.995 ;
    END
  END wd_in_w1[43]
  PIN wd_in_w1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.345 0.070 534.415 ;
    END
  END wd_in_w1[44]
  PIN wd_in_w1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.765 0.070 534.835 ;
    END
  END wd_in_w1[45]
  PIN wd_in_w1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.185 0.070 535.255 ;
    END
  END wd_in_w1[46]
  PIN wd_in_w1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.605 0.070 535.675 ;
    END
  END wd_in_w1[47]
  PIN wd_in_w1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.025 0.070 536.095 ;
    END
  END wd_in_w1[48]
  PIN wd_in_w1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.445 0.070 536.515 ;
    END
  END wd_in_w1[49]
  PIN wd_in_w1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.865 0.070 536.935 ;
    END
  END wd_in_w1[50]
  PIN wd_in_w1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.285 0.070 537.355 ;
    END
  END wd_in_w1[51]
  PIN wd_in_w1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.705 0.070 537.775 ;
    END
  END wd_in_w1[52]
  PIN wd_in_w1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.125 0.070 538.195 ;
    END
  END wd_in_w1[53]
  PIN wd_in_w1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.545 0.070 538.615 ;
    END
  END wd_in_w1[54]
  PIN wd_in_w1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.965 0.070 539.035 ;
    END
  END wd_in_w1[55]
  PIN wd_in_w1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.385 0.070 539.455 ;
    END
  END wd_in_w1[56]
  PIN wd_in_w1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.805 0.070 539.875 ;
    END
  END wd_in_w1[57]
  PIN wd_in_w1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.225 0.070 540.295 ;
    END
  END wd_in_w1[58]
  PIN wd_in_w1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.645 0.070 540.715 ;
    END
  END wd_in_w1[59]
  PIN wd_in_w1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.065 0.070 541.135 ;
    END
  END wd_in_w1[60]
  PIN wd_in_w1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.485 0.070 541.555 ;
    END
  END wd_in_w1[61]
  PIN wd_in_w1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.905 0.070 541.975 ;
    END
  END wd_in_w1[62]
  PIN wd_in_w1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.325 0.070 542.395 ;
    END
  END wd_in_w1[63]
  PIN wd_in_w1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.745 0.070 542.815 ;
    END
  END wd_in_w1[64]
  PIN wd_in_w1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.165 0.070 543.235 ;
    END
  END wd_in_w1[65]
  PIN wd_in_w1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.585 0.070 543.655 ;
    END
  END wd_in_w1[66]
  PIN wd_in_w1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.005 0.070 544.075 ;
    END
  END wd_in_w1[67]
  PIN wd_in_w1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.425 0.070 544.495 ;
    END
  END wd_in_w1[68]
  PIN wd_in_w1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.845 0.070 544.915 ;
    END
  END wd_in_w1[69]
  PIN wd_in_w1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.265 0.070 545.335 ;
    END
  END wd_in_w1[70]
  PIN wd_in_w1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.685 0.070 545.755 ;
    END
  END wd_in_w1[71]
  PIN wd_in_w1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.105 0.070 546.175 ;
    END
  END wd_in_w1[72]
  PIN wd_in_w1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.525 0.070 546.595 ;
    END
  END wd_in_w1[73]
  PIN wd_in_w1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.945 0.070 547.015 ;
    END
  END wd_in_w1[74]
  PIN wd_in_w1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.365 0.070 547.435 ;
    END
  END wd_in_w1[75]
  PIN wd_in_w1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.785 0.070 547.855 ;
    END
  END wd_in_w1[76]
  PIN wd_in_w1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.205 0.070 548.275 ;
    END
  END wd_in_w1[77]
  PIN wd_in_w1[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.625 0.070 548.695 ;
    END
  END wd_in_w1[78]
  PIN wd_in_w1[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.045 0.070 549.115 ;
    END
  END wd_in_w1[79]
  PIN wd_in_w1[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.465 0.070 549.535 ;
    END
  END wd_in_w1[80]
  PIN wd_in_w1[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.885 0.070 549.955 ;
    END
  END wd_in_w1[81]
  PIN wd_in_w1[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.305 0.070 550.375 ;
    END
  END wd_in_w1[82]
  PIN wd_in_w1[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.725 0.070 550.795 ;
    END
  END wd_in_w1[83]
  PIN wd_in_w1[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.145 0.070 551.215 ;
    END
  END wd_in_w1[84]
  PIN wd_in_w1[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.565 0.070 551.635 ;
    END
  END wd_in_w1[85]
  PIN wd_in_w1[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.985 0.070 552.055 ;
    END
  END wd_in_w1[86]
  PIN wd_in_w1[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.405 0.070 552.475 ;
    END
  END wd_in_w1[87]
  PIN wd_in_w1[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.825 0.070 552.895 ;
    END
  END wd_in_w1[88]
  PIN wd_in_w1[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.245 0.070 553.315 ;
    END
  END wd_in_w1[89]
  PIN wd_in_w1[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.665 0.070 553.735 ;
    END
  END wd_in_w1[90]
  PIN wd_in_w1[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.085 0.070 554.155 ;
    END
  END wd_in_w1[91]
  PIN wd_in_w1[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.505 0.070 554.575 ;
    END
  END wd_in_w1[92]
  PIN wd_in_w1[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.925 0.070 554.995 ;
    END
  END wd_in_w1[93]
  PIN wd_in_w1[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.345 0.070 555.415 ;
    END
  END wd_in_w1[94]
  PIN wd_in_w1[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.765 0.070 555.835 ;
    END
  END wd_in_w1[95]
  PIN wd_in_w1[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.185 0.070 556.255 ;
    END
  END wd_in_w1[96]
  PIN wd_in_w1[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.605 0.070 556.675 ;
    END
  END wd_in_w1[97]
  PIN wd_in_w1[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.025 0.070 557.095 ;
    END
  END wd_in_w1[98]
  PIN wd_in_w1[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.445 0.070 557.515 ;
    END
  END wd_in_w1[99]
  PIN wd_in_w1[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.865 0.070 557.935 ;
    END
  END wd_in_w1[100]
  PIN wd_in_w1[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.285 0.070 558.355 ;
    END
  END wd_in_w1[101]
  PIN wd_in_w1[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.705 0.070 558.775 ;
    END
  END wd_in_w1[102]
  PIN wd_in_w1[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.125 0.070 559.195 ;
    END
  END wd_in_w1[103]
  PIN wd_in_w1[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.545 0.070 559.615 ;
    END
  END wd_in_w1[104]
  PIN wd_in_w1[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.965 0.070 560.035 ;
    END
  END wd_in_w1[105]
  PIN wd_in_w1[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.385 0.070 560.455 ;
    END
  END wd_in_w1[106]
  PIN wd_in_w1[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.805 0.070 560.875 ;
    END
  END wd_in_w1[107]
  PIN wd_in_w1[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.225 0.070 561.295 ;
    END
  END wd_in_w1[108]
  PIN wd_in_w1[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.645 0.070 561.715 ;
    END
  END wd_in_w1[109]
  PIN wd_in_w1[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.065 0.070 562.135 ;
    END
  END wd_in_w1[110]
  PIN wd_in_w1[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.485 0.070 562.555 ;
    END
  END wd_in_w1[111]
  PIN wd_in_w1[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.905 0.070 562.975 ;
    END
  END wd_in_w1[112]
  PIN wd_in_w1[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.325 0.070 563.395 ;
    END
  END wd_in_w1[113]
  PIN wd_in_w1[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.745 0.070 563.815 ;
    END
  END wd_in_w1[114]
  PIN wd_in_w1[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.165 0.070 564.235 ;
    END
  END wd_in_w1[115]
  PIN wd_in_w1[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.585 0.070 564.655 ;
    END
  END wd_in_w1[116]
  PIN wd_in_w1[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.005 0.070 565.075 ;
    END
  END wd_in_w1[117]
  PIN wd_in_w1[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.425 0.070 565.495 ;
    END
  END wd_in_w1[118]
  PIN wd_in_w1[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.845 0.070 565.915 ;
    END
  END wd_in_w1[119]
  PIN wd_in_w1[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.265 0.070 566.335 ;
    END
  END wd_in_w1[120]
  PIN wd_in_w1[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.685 0.070 566.755 ;
    END
  END wd_in_w1[121]
  PIN wd_in_w1[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.105 0.070 567.175 ;
    END
  END wd_in_w1[122]
  PIN wd_in_w1[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.525 0.070 567.595 ;
    END
  END wd_in_w1[123]
  PIN wd_in_w1[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.945 0.070 568.015 ;
    END
  END wd_in_w1[124]
  PIN wd_in_w1[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.365 0.070 568.435 ;
    END
  END wd_in_w1[125]
  PIN wd_in_w1[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.785 0.070 568.855 ;
    END
  END wd_in_w1[126]
  PIN wd_in_w1[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.205 0.070 569.275 ;
    END
  END wd_in_w1[127]
  PIN wd_in_w1[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.625 0.070 569.695 ;
    END
  END wd_in_w1[128]
  PIN wd_in_w1[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.045 0.070 570.115 ;
    END
  END wd_in_w1[129]
  PIN wd_in_w1[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.465 0.070 570.535 ;
    END
  END wd_in_w1[130]
  PIN wd_in_w1[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.885 0.070 570.955 ;
    END
  END wd_in_w1[131]
  PIN wd_in_w1[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.305 0.070 571.375 ;
    END
  END wd_in_w1[132]
  PIN wd_in_w1[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.725 0.070 571.795 ;
    END
  END wd_in_w1[133]
  PIN wd_in_w1[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.145 0.070 572.215 ;
    END
  END wd_in_w1[134]
  PIN wd_in_w1[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.565 0.070 572.635 ;
    END
  END wd_in_w1[135]
  PIN wd_in_w1[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.985 0.070 573.055 ;
    END
  END wd_in_w1[136]
  PIN wd_in_w1[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.405 0.070 573.475 ;
    END
  END wd_in_w1[137]
  PIN wd_in_w1[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.825 0.070 573.895 ;
    END
  END wd_in_w1[138]
  PIN wd_in_w1[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.245 0.070 574.315 ;
    END
  END wd_in_w1[139]
  PIN wd_in_w1[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.665 0.070 574.735 ;
    END
  END wd_in_w1[140]
  PIN wd_in_w1[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.085 0.070 575.155 ;
    END
  END wd_in_w1[141]
  PIN wd_in_w1[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.505 0.070 575.575 ;
    END
  END wd_in_w1[142]
  PIN wd_in_w1[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.925 0.070 575.995 ;
    END
  END wd_in_w1[143]
  PIN wd_in_w1[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 576.345 0.070 576.415 ;
    END
  END wd_in_w1[144]
  PIN wd_in_w1[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 576.765 0.070 576.835 ;
    END
  END wd_in_w1[145]
  PIN wd_in_w1[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.185 0.070 577.255 ;
    END
  END wd_in_w1[146]
  PIN wd_in_w1[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.605 0.070 577.675 ;
    END
  END wd_in_w1[147]
  PIN wd_in_w1[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.025 0.070 578.095 ;
    END
  END wd_in_w1[148]
  PIN wd_in_w1[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.445 0.070 578.515 ;
    END
  END wd_in_w1[149]
  PIN wd_in_w1[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.865 0.070 578.935 ;
    END
  END wd_in_w1[150]
  PIN wd_in_w1[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.285 0.070 579.355 ;
    END
  END wd_in_w1[151]
  PIN wd_in_w1[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.705 0.070 579.775 ;
    END
  END wd_in_w1[152]
  PIN wd_in_w1[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.125 0.070 580.195 ;
    END
  END wd_in_w1[153]
  PIN wd_in_w1[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.545 0.070 580.615 ;
    END
  END wd_in_w1[154]
  PIN wd_in_w1[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.965 0.070 581.035 ;
    END
  END wd_in_w1[155]
  PIN wd_in_w1[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 581.385 0.070 581.455 ;
    END
  END wd_in_w1[156]
  PIN wd_in_w1[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 581.805 0.070 581.875 ;
    END
  END wd_in_w1[157]
  PIN wd_in_w1[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.225 0.070 582.295 ;
    END
  END wd_in_w1[158]
  PIN wd_in_w1[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.645 0.070 582.715 ;
    END
  END wd_in_w1[159]
  PIN wd_in_w1[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.065 0.070 583.135 ;
    END
  END wd_in_w1[160]
  PIN wd_in_w1[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.485 0.070 583.555 ;
    END
  END wd_in_w1[161]
  PIN wd_in_w1[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.905 0.070 583.975 ;
    END
  END wd_in_w1[162]
  PIN wd_in_w1[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.325 0.070 584.395 ;
    END
  END wd_in_w1[163]
  PIN wd_in_w1[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.745 0.070 584.815 ;
    END
  END wd_in_w1[164]
  PIN wd_in_w1[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 585.165 0.070 585.235 ;
    END
  END wd_in_w1[165]
  PIN wd_in_w1[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 585.585 0.070 585.655 ;
    END
  END wd_in_w1[166]
  PIN wd_in_w1[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.005 0.070 586.075 ;
    END
  END wd_in_w1[167]
  PIN wd_in_w1[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.425 0.070 586.495 ;
    END
  END wd_in_w1[168]
  PIN wd_in_w1[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.845 0.070 586.915 ;
    END
  END wd_in_w1[169]
  PIN wd_in_w1[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.265 0.070 587.335 ;
    END
  END wd_in_w1[170]
  PIN wd_in_w1[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.685 0.070 587.755 ;
    END
  END wd_in_w1[171]
  PIN wd_in_w1[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.105 0.070 588.175 ;
    END
  END wd_in_w1[172]
  PIN wd_in_w1[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.525 0.070 588.595 ;
    END
  END wd_in_w1[173]
  PIN wd_in_w1[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.945 0.070 589.015 ;
    END
  END wd_in_w1[174]
  PIN wd_in_w1[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.365 0.070 589.435 ;
    END
  END wd_in_w1[175]
  PIN wd_in_w1[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.785 0.070 589.855 ;
    END
  END wd_in_w1[176]
  PIN wd_in_w1[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 590.205 0.070 590.275 ;
    END
  END wd_in_w1[177]
  PIN wd_in_w1[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 590.625 0.070 590.695 ;
    END
  END wd_in_w1[178]
  PIN wd_in_w1[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.045 0.070 591.115 ;
    END
  END wd_in_w1[179]
  PIN wd_in_w1[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.465 0.070 591.535 ;
    END
  END wd_in_w1[180]
  PIN wd_in_w1[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.885 0.070 591.955 ;
    END
  END wd_in_w1[181]
  PIN wd_in_w1[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.305 0.070 592.375 ;
    END
  END wd_in_w1[182]
  PIN wd_in_w1[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.725 0.070 592.795 ;
    END
  END wd_in_w1[183]
  PIN wd_in_w1[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.145 0.070 593.215 ;
    END
  END wd_in_w1[184]
  PIN wd_in_w1[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.565 0.070 593.635 ;
    END
  END wd_in_w1[185]
  PIN wd_in_w1[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.985 0.070 594.055 ;
    END
  END wd_in_w1[186]
  PIN wd_in_w1[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.405 0.070 594.475 ;
    END
  END wd_in_w1[187]
  PIN wd_in_w1[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.825 0.070 594.895 ;
    END
  END wd_in_w1[188]
  PIN wd_in_w1[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.245 0.070 595.315 ;
    END
  END wd_in_w1[189]
  PIN wd_in_w1[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.665 0.070 595.735 ;
    END
  END wd_in_w1[190]
  PIN wd_in_w1[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.085 0.070 596.155 ;
    END
  END wd_in_w1[191]
  PIN wd_in_w1[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.505 0.070 596.575 ;
    END
  END wd_in_w1[192]
  PIN wd_in_w1[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.925 0.070 596.995 ;
    END
  END wd_in_w1[193]
  PIN wd_in_w1[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.345 0.070 597.415 ;
    END
  END wd_in_w1[194]
  PIN wd_in_w1[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.765 0.070 597.835 ;
    END
  END wd_in_w1[195]
  PIN wd_in_w1[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.185 0.070 598.255 ;
    END
  END wd_in_w1[196]
  PIN wd_in_w1[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.605 0.070 598.675 ;
    END
  END wd_in_w1[197]
  PIN wd_in_w1[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.025 0.070 599.095 ;
    END
  END wd_in_w1[198]
  PIN wd_in_w1[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.445 0.070 599.515 ;
    END
  END wd_in_w1[199]
  PIN wd_in_w1[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.865 0.070 599.935 ;
    END
  END wd_in_w1[200]
  PIN wd_in_w1[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.285 0.070 600.355 ;
    END
  END wd_in_w1[201]
  PIN wd_in_w1[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.705 0.070 600.775 ;
    END
  END wd_in_w1[202]
  PIN wd_in_w1[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.125 0.070 601.195 ;
    END
  END wd_in_w1[203]
  PIN wd_in_w1[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.545 0.070 601.615 ;
    END
  END wd_in_w1[204]
  PIN wd_in_w1[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.965 0.070 602.035 ;
    END
  END wd_in_w1[205]
  PIN wd_in_w1[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.385 0.070 602.455 ;
    END
  END wd_in_w1[206]
  PIN wd_in_w1[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.805 0.070 602.875 ;
    END
  END wd_in_w1[207]
  PIN wd_in_w1[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.225 0.070 603.295 ;
    END
  END wd_in_w1[208]
  PIN wd_in_w1[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.645 0.070 603.715 ;
    END
  END wd_in_w1[209]
  PIN wd_in_w1[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.065 0.070 604.135 ;
    END
  END wd_in_w1[210]
  PIN wd_in_w1[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.485 0.070 604.555 ;
    END
  END wd_in_w1[211]
  PIN wd_in_w1[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.905 0.070 604.975 ;
    END
  END wd_in_w1[212]
  PIN wd_in_w1[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.325 0.070 605.395 ;
    END
  END wd_in_w1[213]
  PIN wd_in_w1[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.745 0.070 605.815 ;
    END
  END wd_in_w1[214]
  PIN wd_in_w1[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.165 0.070 606.235 ;
    END
  END wd_in_w1[215]
  PIN wd_in_w1[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.585 0.070 606.655 ;
    END
  END wd_in_w1[216]
  PIN wd_in_w1[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.005 0.070 607.075 ;
    END
  END wd_in_w1[217]
  PIN wd_in_w1[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.425 0.070 607.495 ;
    END
  END wd_in_w1[218]
  PIN wd_in_w1[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.845 0.070 607.915 ;
    END
  END wd_in_w1[219]
  PIN wd_in_w1[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.265 0.070 608.335 ;
    END
  END wd_in_w1[220]
  PIN wd_in_w1[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.685 0.070 608.755 ;
    END
  END wd_in_w1[221]
  PIN wd_in_w1[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.105 0.070 609.175 ;
    END
  END wd_in_w1[222]
  PIN wd_in_w1[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.525 0.070 609.595 ;
    END
  END wd_in_w1[223]
  PIN wd_in_w1[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.945 0.070 610.015 ;
    END
  END wd_in_w1[224]
  PIN wd_in_w1[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.365 0.070 610.435 ;
    END
  END wd_in_w1[225]
  PIN wd_in_w1[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.785 0.070 610.855 ;
    END
  END wd_in_w1[226]
  PIN wd_in_w1[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.205 0.070 611.275 ;
    END
  END wd_in_w1[227]
  PIN wd_in_w1[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.625 0.070 611.695 ;
    END
  END wd_in_w1[228]
  PIN wd_in_w1[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.045 0.070 612.115 ;
    END
  END wd_in_w1[229]
  PIN wd_in_w1[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.465 0.070 612.535 ;
    END
  END wd_in_w1[230]
  PIN wd_in_w1[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.885 0.070 612.955 ;
    END
  END wd_in_w1[231]
  PIN wd_in_w1[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 613.305 0.070 613.375 ;
    END
  END wd_in_w1[232]
  PIN wd_in_w1[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 613.725 0.070 613.795 ;
    END
  END wd_in_w1[233]
  PIN wd_in_w1[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.145 0.070 614.215 ;
    END
  END wd_in_w1[234]
  PIN wd_in_w1[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.565 0.070 614.635 ;
    END
  END wd_in_w1[235]
  PIN wd_in_w1[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.985 0.070 615.055 ;
    END
  END wd_in_w1[236]
  PIN wd_in_w1[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.405 0.070 615.475 ;
    END
  END wd_in_w1[237]
  PIN wd_in_w1[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.825 0.070 615.895 ;
    END
  END wd_in_w1[238]
  PIN wd_in_w1[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.245 0.070 616.315 ;
    END
  END wd_in_w1[239]
  PIN wd_in_w1[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.665 0.070 616.735 ;
    END
  END wd_in_w1[240]
  PIN wd_in_w1[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.085 0.070 617.155 ;
    END
  END wd_in_w1[241]
  PIN wd_in_w1[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.505 0.070 617.575 ;
    END
  END wd_in_w1[242]
  PIN wd_in_w1[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.925 0.070 617.995 ;
    END
  END wd_in_w1[243]
  PIN wd_in_w1[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.345 0.070 618.415 ;
    END
  END wd_in_w1[244]
  PIN wd_in_w1[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.765 0.070 618.835 ;
    END
  END wd_in_w1[245]
  PIN wd_in_w1[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.185 0.070 619.255 ;
    END
  END wd_in_w1[246]
  PIN wd_in_w1[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.605 0.070 619.675 ;
    END
  END wd_in_w1[247]
  PIN wd_in_w1[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.025 0.070 620.095 ;
    END
  END wd_in_w1[248]
  PIN wd_in_w1[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.445 0.070 620.515 ;
    END
  END wd_in_w1[249]
  PIN wd_in_w1[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.865 0.070 620.935 ;
    END
  END wd_in_w1[250]
  PIN wd_in_w1[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.285 0.070 621.355 ;
    END
  END wd_in_w1[251]
  PIN wd_in_w1[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.705 0.070 621.775 ;
    END
  END wd_in_w1[252]
  PIN wd_in_w1[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.125 0.070 622.195 ;
    END
  END wd_in_w1[253]
  PIN wd_in_w1[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.545 0.070 622.615 ;
    END
  END wd_in_w1[254]
  PIN wd_in_w1[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.965 0.070 623.035 ;
    END
  END wd_in_w1[255]
  PIN wd_in_w1[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.385 0.070 623.455 ;
    END
  END wd_in_w1[256]
  PIN wd_in_w1[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.805 0.070 623.875 ;
    END
  END wd_in_w1[257]
  PIN wd_in_w1[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.225 0.070 624.295 ;
    END
  END wd_in_w1[258]
  PIN wd_in_w1[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.645 0.070 624.715 ;
    END
  END wd_in_w1[259]
  PIN wd_in_w1[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.065 0.070 625.135 ;
    END
  END wd_in_w1[260]
  PIN wd_in_w1[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.485 0.070 625.555 ;
    END
  END wd_in_w1[261]
  PIN wd_in_w1[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.905 0.070 625.975 ;
    END
  END wd_in_w1[262]
  PIN wd_in_w1[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.325 0.070 626.395 ;
    END
  END wd_in_w1[263]
  PIN wd_in_w1[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.745 0.070 626.815 ;
    END
  END wd_in_w1[264]
  PIN wd_in_w1[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 627.165 0.070 627.235 ;
    END
  END wd_in_w1[265]
  PIN wd_in_w1[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 627.585 0.070 627.655 ;
    END
  END wd_in_w1[266]
  PIN wd_in_w1[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.005 0.070 628.075 ;
    END
  END wd_in_w1[267]
  PIN wd_in_w1[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.425 0.070 628.495 ;
    END
  END wd_in_w1[268]
  PIN wd_in_w1[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.845 0.070 628.915 ;
    END
  END wd_in_w1[269]
  PIN wd_in_w1[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 629.265 0.070 629.335 ;
    END
  END wd_in_w1[270]
  PIN wd_in_w1[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 629.685 0.070 629.755 ;
    END
  END wd_in_w1[271]
  PIN wd_in_w1[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 630.105 0.070 630.175 ;
    END
  END wd_in_w1[272]
  PIN wd_in_w1[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 630.525 0.070 630.595 ;
    END
  END wd_in_w1[273]
  PIN wd_in_w1[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 630.945 0.070 631.015 ;
    END
  END wd_in_w1[274]
  PIN wd_in_w1[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.365 0.070 631.435 ;
    END
  END wd_in_w1[275]
  PIN wd_in_w1[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.785 0.070 631.855 ;
    END
  END wd_in_w1[276]
  PIN wd_in_w1[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 632.205 0.070 632.275 ;
    END
  END wd_in_w1[277]
  PIN wd_in_w1[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 632.625 0.070 632.695 ;
    END
  END wd_in_w1[278]
  PIN wd_in_w1[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.045 0.070 633.115 ;
    END
  END wd_in_w1[279]
  PIN wd_in_w1[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.465 0.070 633.535 ;
    END
  END wd_in_w1[280]
  PIN wd_in_w1[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.885 0.070 633.955 ;
    END
  END wd_in_w1[281]
  PIN wd_in_w1[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 634.305 0.070 634.375 ;
    END
  END wd_in_w1[282]
  PIN wd_in_w1[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 634.725 0.070 634.795 ;
    END
  END wd_in_w1[283]
  PIN wd_in_w1[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.145 0.070 635.215 ;
    END
  END wd_in_w1[284]
  PIN wd_in_w1[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.565 0.070 635.635 ;
    END
  END wd_in_w1[285]
  PIN wd_in_w1[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.985 0.070 636.055 ;
    END
  END wd_in_w1[286]
  PIN wd_in_w1[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.405 0.070 636.475 ;
    END
  END wd_in_w1[287]
  PIN wd_in_w1[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.825 0.070 636.895 ;
    END
  END wd_in_w1[288]
  PIN wd_in_w1[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 637.245 0.070 637.315 ;
    END
  END wd_in_w1[289]
  PIN wd_in_w1[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 637.665 0.070 637.735 ;
    END
  END wd_in_w1[290]
  PIN wd_in_w1[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.085 0.070 638.155 ;
    END
  END wd_in_w1[291]
  PIN wd_in_w1[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.505 0.070 638.575 ;
    END
  END wd_in_w1[292]
  PIN wd_in_w1[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.925 0.070 638.995 ;
    END
  END wd_in_w1[293]
  PIN wd_in_w1[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 639.345 0.070 639.415 ;
    END
  END wd_in_w1[294]
  PIN wd_in_w1[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 639.765 0.070 639.835 ;
    END
  END wd_in_w1[295]
  PIN wd_in_w1[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 640.185 0.070 640.255 ;
    END
  END wd_in_w1[296]
  PIN wd_in_w1[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 640.605 0.070 640.675 ;
    END
  END wd_in_w1[297]
  PIN wd_in_w1[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.025 0.070 641.095 ;
    END
  END wd_in_w1[298]
  PIN wd_in_w1[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.445 0.070 641.515 ;
    END
  END wd_in_w1[299]
  PIN wd_in_w1[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.865 0.070 641.935 ;
    END
  END wd_in_w1[300]
  PIN wd_in_w1[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.285 0.070 642.355 ;
    END
  END wd_in_w1[301]
  PIN wd_in_w1[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.705 0.070 642.775 ;
    END
  END wd_in_w1[302]
  PIN wd_in_w1[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 643.125 0.070 643.195 ;
    END
  END wd_in_w1[303]
  PIN wd_in_w1[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 643.545 0.070 643.615 ;
    END
  END wd_in_w1[304]
  PIN wd_in_w1[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 643.965 0.070 644.035 ;
    END
  END wd_in_w1[305]
  PIN wd_in_w1[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 644.385 0.070 644.455 ;
    END
  END wd_in_w1[306]
  PIN wd_in_w1[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 644.805 0.070 644.875 ;
    END
  END wd_in_w1[307]
  PIN wd_in_w1[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 645.225 0.070 645.295 ;
    END
  END wd_in_w1[308]
  PIN wd_in_w1[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 645.645 0.070 645.715 ;
    END
  END wd_in_w1[309]
  PIN wd_in_w1[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.065 0.070 646.135 ;
    END
  END wd_in_w1[310]
  PIN wd_in_w1[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.485 0.070 646.555 ;
    END
  END wd_in_w1[311]
  PIN wd_in_w1[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.905 0.070 646.975 ;
    END
  END wd_in_w1[312]
  PIN wd_in_w1[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.325 0.070 647.395 ;
    END
  END wd_in_w1[313]
  PIN wd_in_w1[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.745 0.070 647.815 ;
    END
  END wd_in_w1[314]
  PIN wd_in_w1[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 648.165 0.070 648.235 ;
    END
  END wd_in_w1[315]
  PIN wd_in_w1[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 648.585 0.070 648.655 ;
    END
  END wd_in_w1[316]
  PIN wd_in_w1[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.005 0.070 649.075 ;
    END
  END wd_in_w1[317]
  PIN wd_in_w1[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.425 0.070 649.495 ;
    END
  END wd_in_w1[318]
  PIN wd_in_w1[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.845 0.070 649.915 ;
    END
  END wd_in_w1[319]
  PIN wd_in_w1[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 650.265 0.070 650.335 ;
    END
  END wd_in_w1[320]
  PIN wd_in_w1[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 650.685 0.070 650.755 ;
    END
  END wd_in_w1[321]
  PIN wd_in_w1[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 651.105 0.070 651.175 ;
    END
  END wd_in_w1[322]
  PIN wd_in_w1[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 651.525 0.070 651.595 ;
    END
  END wd_in_w1[323]
  PIN wd_in_w1[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 651.945 0.070 652.015 ;
    END
  END wd_in_w1[324]
  PIN wd_in_w1[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.365 0.070 652.435 ;
    END
  END wd_in_w1[325]
  PIN wd_in_w1[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.785 0.070 652.855 ;
    END
  END wd_in_w1[326]
  PIN wd_in_w1[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 653.205 0.070 653.275 ;
    END
  END wd_in_w1[327]
  PIN wd_in_w1[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 653.625 0.070 653.695 ;
    END
  END wd_in_w1[328]
  PIN wd_in_w1[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.045 0.070 654.115 ;
    END
  END wd_in_w1[329]
  PIN wd_in_w1[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.465 0.070 654.535 ;
    END
  END wd_in_w1[330]
  PIN wd_in_w1[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.885 0.070 654.955 ;
    END
  END wd_in_w1[331]
  PIN wd_in_w1[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 655.305 0.070 655.375 ;
    END
  END wd_in_w1[332]
  PIN wd_in_w1[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 655.725 0.070 655.795 ;
    END
  END wd_in_w1[333]
  PIN wd_in_w1[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.145 0.070 656.215 ;
    END
  END wd_in_w1[334]
  PIN wd_in_w1[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.565 0.070 656.635 ;
    END
  END wd_in_w1[335]
  PIN wd_in_w1[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.985 0.070 657.055 ;
    END
  END wd_in_w1[336]
  PIN wd_in_w1[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.405 0.070 657.475 ;
    END
  END wd_in_w1[337]
  PIN wd_in_w1[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.825 0.070 657.895 ;
    END
  END wd_in_w1[338]
  PIN wd_in_w1[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.245 0.070 658.315 ;
    END
  END wd_in_w1[339]
  PIN wd_in_w1[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.665 0.070 658.735 ;
    END
  END wd_in_w1[340]
  PIN wd_in_w1[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.085 0.070 659.155 ;
    END
  END wd_in_w1[341]
  PIN wd_in_w1[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.505 0.070 659.575 ;
    END
  END wd_in_w1[342]
  PIN wd_in_w1[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.925 0.070 659.995 ;
    END
  END wd_in_w1[343]
  PIN wd_in_w1[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.345 0.070 660.415 ;
    END
  END wd_in_w1[344]
  PIN wd_in_w1[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.765 0.070 660.835 ;
    END
  END wd_in_w1[345]
  PIN wd_in_w1[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.185 0.070 661.255 ;
    END
  END wd_in_w1[346]
  PIN wd_in_w1[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.605 0.070 661.675 ;
    END
  END wd_in_w1[347]
  PIN wd_in_w1[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.025 0.070 662.095 ;
    END
  END wd_in_w1[348]
  PIN wd_in_w1[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.445 0.070 662.515 ;
    END
  END wd_in_w1[349]
  PIN wd_in_w1[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.865 0.070 662.935 ;
    END
  END wd_in_w1[350]
  PIN wd_in_w1[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.285 0.070 663.355 ;
    END
  END wd_in_w1[351]
  PIN wd_in_w1[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.705 0.070 663.775 ;
    END
  END wd_in_w1[352]
  PIN wd_in_w1[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.125 0.070 664.195 ;
    END
  END wd_in_w1[353]
  PIN wd_in_w1[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.545 0.070 664.615 ;
    END
  END wd_in_w1[354]
  PIN wd_in_w1[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.965 0.070 665.035 ;
    END
  END wd_in_w1[355]
  PIN wd_in_w1[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.385 0.070 665.455 ;
    END
  END wd_in_w1[356]
  PIN wd_in_w1[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.805 0.070 665.875 ;
    END
  END wd_in_w1[357]
  PIN wd_in_w1[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.225 0.070 666.295 ;
    END
  END wd_in_w1[358]
  PIN wd_in_w1[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.645 0.070 666.715 ;
    END
  END wd_in_w1[359]
  PIN wd_in_w1[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.065 0.070 667.135 ;
    END
  END wd_in_w1[360]
  PIN wd_in_w1[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.485 0.070 667.555 ;
    END
  END wd_in_w1[361]
  PIN wd_in_w1[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.905 0.070 667.975 ;
    END
  END wd_in_w1[362]
  PIN wd_in_w1[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.325 0.070 668.395 ;
    END
  END wd_in_w1[363]
  PIN wd_in_w1[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.745 0.070 668.815 ;
    END
  END wd_in_w1[364]
  PIN wd_in_w1[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.165 0.070 669.235 ;
    END
  END wd_in_w1[365]
  PIN wd_in_w1[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.585 0.070 669.655 ;
    END
  END wd_in_w1[366]
  PIN wd_in_w1[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.005 0.070 670.075 ;
    END
  END wd_in_w1[367]
  PIN wd_in_w1[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.425 0.070 670.495 ;
    END
  END wd_in_w1[368]
  PIN wd_in_w1[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.845 0.070 670.915 ;
    END
  END wd_in_w1[369]
  PIN wd_in_w1[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.265 0.070 671.335 ;
    END
  END wd_in_w1[370]
  PIN wd_in_w1[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.685 0.070 671.755 ;
    END
  END wd_in_w1[371]
  PIN wd_in_w1[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.105 0.070 672.175 ;
    END
  END wd_in_w1[372]
  PIN wd_in_w1[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.525 0.070 672.595 ;
    END
  END wd_in_w1[373]
  PIN wd_in_w1[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.945 0.070 673.015 ;
    END
  END wd_in_w1[374]
  PIN wd_in_w1[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.365 0.070 673.435 ;
    END
  END wd_in_w1[375]
  PIN wd_in_w1[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.785 0.070 673.855 ;
    END
  END wd_in_w1[376]
  PIN wd_in_w1[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.205 0.070 674.275 ;
    END
  END wd_in_w1[377]
  PIN wd_in_w1[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.625 0.070 674.695 ;
    END
  END wd_in_w1[378]
  PIN wd_in_w1[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.045 0.070 675.115 ;
    END
  END wd_in_w1[379]
  PIN wd_in_w1[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.465 0.070 675.535 ;
    END
  END wd_in_w1[380]
  PIN wd_in_w1[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.885 0.070 675.955 ;
    END
  END wd_in_w1[381]
  PIN wd_in_w1[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 676.305 0.070 676.375 ;
    END
  END wd_in_w1[382]
  PIN wd_in_w1[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 676.725 0.070 676.795 ;
    END
  END wd_in_w1[383]
  PIN wd_in_w1[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.145 0.070 677.215 ;
    END
  END wd_in_w1[384]
  PIN wd_in_w1[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.565 0.070 677.635 ;
    END
  END wd_in_w1[385]
  PIN wd_in_w1[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.985 0.070 678.055 ;
    END
  END wd_in_w1[386]
  PIN wd_in_w1[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.405 0.070 678.475 ;
    END
  END wd_in_w1[387]
  PIN wd_in_w1[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.825 0.070 678.895 ;
    END
  END wd_in_w1[388]
  PIN wd_in_w1[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.245 0.070 679.315 ;
    END
  END wd_in_w1[389]
  PIN wd_in_w1[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.665 0.070 679.735 ;
    END
  END wd_in_w1[390]
  PIN wd_in_w1[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.085 0.070 680.155 ;
    END
  END wd_in_w1[391]
  PIN wd_in_w1[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.505 0.070 680.575 ;
    END
  END wd_in_w1[392]
  PIN wd_in_w1[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.925 0.070 680.995 ;
    END
  END wd_in_w1[393]
  PIN wd_in_w1[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.345 0.070 681.415 ;
    END
  END wd_in_w1[394]
  PIN wd_in_w1[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.765 0.070 681.835 ;
    END
  END wd_in_w1[395]
  PIN wd_in_w1[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.185 0.070 682.255 ;
    END
  END wd_in_w1[396]
  PIN wd_in_w1[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.605 0.070 682.675 ;
    END
  END wd_in_w1[397]
  PIN wd_in_w1[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.025 0.070 683.095 ;
    END
  END wd_in_w1[398]
  PIN wd_in_w1[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.445 0.070 683.515 ;
    END
  END wd_in_w1[399]
  PIN wd_in_w1[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.865 0.070 683.935 ;
    END
  END wd_in_w1[400]
  PIN wd_in_w1[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.285 0.070 684.355 ;
    END
  END wd_in_w1[401]
  PIN wd_in_w1[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.705 0.070 684.775 ;
    END
  END wd_in_w1[402]
  PIN wd_in_w1[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.125 0.070 685.195 ;
    END
  END wd_in_w1[403]
  PIN wd_in_w1[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.545 0.070 685.615 ;
    END
  END wd_in_w1[404]
  PIN wd_in_w1[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.965 0.070 686.035 ;
    END
  END wd_in_w1[405]
  PIN wd_in_w1[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 686.385 0.070 686.455 ;
    END
  END wd_in_w1[406]
  PIN wd_in_w1[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 686.805 0.070 686.875 ;
    END
  END wd_in_w1[407]
  PIN wd_in_w1[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.225 0.070 687.295 ;
    END
  END wd_in_w1[408]
  PIN wd_in_w1[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.645 0.070 687.715 ;
    END
  END wd_in_w1[409]
  PIN wd_in_w1[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.065 0.070 688.135 ;
    END
  END wd_in_w1[410]
  PIN wd_in_w1[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.485 0.070 688.555 ;
    END
  END wd_in_w1[411]
  PIN wd_in_w1[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.905 0.070 688.975 ;
    END
  END wd_in_w1[412]
  PIN wd_in_w1[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.325 0.070 689.395 ;
    END
  END wd_in_w1[413]
  PIN wd_in_w1[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.745 0.070 689.815 ;
    END
  END wd_in_w1[414]
  PIN wd_in_w1[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 690.165 0.070 690.235 ;
    END
  END wd_in_w1[415]
  PIN wd_in_w1[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 690.585 0.070 690.655 ;
    END
  END wd_in_w1[416]
  PIN wd_in_w1[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.005 0.070 691.075 ;
    END
  END wd_in_w1[417]
  PIN wd_in_w1[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.425 0.070 691.495 ;
    END
  END wd_in_w1[418]
  PIN wd_in_w1[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.845 0.070 691.915 ;
    END
  END wd_in_w1[419]
  PIN wd_in_w1[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.265 0.070 692.335 ;
    END
  END wd_in_w1[420]
  PIN wd_in_w1[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.685 0.070 692.755 ;
    END
  END wd_in_w1[421]
  PIN wd_in_w1[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.105 0.070 693.175 ;
    END
  END wd_in_w1[422]
  PIN wd_in_w1[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.525 0.070 693.595 ;
    END
  END wd_in_w1[423]
  PIN wd_in_w1[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.945 0.070 694.015 ;
    END
  END wd_in_w1[424]
  PIN wd_in_w1[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.365 0.070 694.435 ;
    END
  END wd_in_w1[425]
  PIN wd_in_w1[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.785 0.070 694.855 ;
    END
  END wd_in_w1[426]
  PIN wd_in_w1[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 695.205 0.070 695.275 ;
    END
  END wd_in_w1[427]
  PIN wd_in_w1[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 695.625 0.070 695.695 ;
    END
  END wd_in_w1[428]
  PIN wd_in_w1[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.045 0.070 696.115 ;
    END
  END wd_in_w1[429]
  PIN wd_in_w1[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.465 0.070 696.535 ;
    END
  END wd_in_w1[430]
  PIN wd_in_w1[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.885 0.070 696.955 ;
    END
  END wd_in_w1[431]
  PIN wd_in_w1[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 697.305 0.070 697.375 ;
    END
  END wd_in_w1[432]
  PIN wd_in_w1[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 697.725 0.070 697.795 ;
    END
  END wd_in_w1[433]
  PIN wd_in_w1[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.145 0.070 698.215 ;
    END
  END wd_in_w1[434]
  PIN wd_in_w1[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.565 0.070 698.635 ;
    END
  END wd_in_w1[435]
  PIN wd_in_w1[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.985 0.070 699.055 ;
    END
  END wd_in_w1[436]
  PIN wd_in_w1[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 699.405 0.070 699.475 ;
    END
  END wd_in_w1[437]
  PIN wd_in_w1[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 699.825 0.070 699.895 ;
    END
  END wd_in_w1[438]
  PIN wd_in_w1[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 700.245 0.070 700.315 ;
    END
  END wd_in_w1[439]
  PIN wd_in_w1[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 700.665 0.070 700.735 ;
    END
  END wd_in_w1[440]
  PIN wd_in_w1[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.085 0.070 701.155 ;
    END
  END wd_in_w1[441]
  PIN wd_in_w1[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.505 0.070 701.575 ;
    END
  END wd_in_w1[442]
  PIN wd_in_w1[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.925 0.070 701.995 ;
    END
  END wd_in_w1[443]
  PIN wd_in_w1[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.345 0.070 702.415 ;
    END
  END wd_in_w1[444]
  PIN wd_in_w1[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.765 0.070 702.835 ;
    END
  END wd_in_w1[445]
  PIN wd_in_w1[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.185 0.070 703.255 ;
    END
  END wd_in_w1[446]
  PIN wd_in_w1[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.605 0.070 703.675 ;
    END
  END wd_in_w1[447]
  PIN wd_in_w1[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.025 0.070 704.095 ;
    END
  END wd_in_w1[448]
  PIN wd_in_w1[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.445 0.070 704.515 ;
    END
  END wd_in_w1[449]
  PIN wd_in_w1[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.865 0.070 704.935 ;
    END
  END wd_in_w1[450]
  PIN wd_in_w1[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.285 0.070 705.355 ;
    END
  END wd_in_w1[451]
  PIN wd_in_w1[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.705 0.070 705.775 ;
    END
  END wd_in_w1[452]
  PIN wd_in_w1[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.125 0.070 706.195 ;
    END
  END wd_in_w1[453]
  PIN wd_in_w1[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.545 0.070 706.615 ;
    END
  END wd_in_w1[454]
  PIN wd_in_w1[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.965 0.070 707.035 ;
    END
  END wd_in_w1[455]
  PIN wd_in_w1[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.385 0.070 707.455 ;
    END
  END wd_in_w1[456]
  PIN wd_in_w1[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.805 0.070 707.875 ;
    END
  END wd_in_w1[457]
  PIN wd_in_w1[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.225 0.070 708.295 ;
    END
  END wd_in_w1[458]
  PIN wd_in_w1[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.645 0.070 708.715 ;
    END
  END wd_in_w1[459]
  PIN wd_in_w1[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.065 0.070 709.135 ;
    END
  END wd_in_w1[460]
  PIN wd_in_w1[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.485 0.070 709.555 ;
    END
  END wd_in_w1[461]
  PIN wd_in_w1[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.905 0.070 709.975 ;
    END
  END wd_in_w1[462]
  PIN wd_in_w1[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.325 0.070 710.395 ;
    END
  END wd_in_w1[463]
  PIN wd_in_w1[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.745 0.070 710.815 ;
    END
  END wd_in_w1[464]
  PIN wd_in_w1[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 711.165 0.070 711.235 ;
    END
  END wd_in_w1[465]
  PIN wd_in_w1[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 711.585 0.070 711.655 ;
    END
  END wd_in_w1[466]
  PIN wd_in_w1[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.005 0.070 712.075 ;
    END
  END wd_in_w1[467]
  PIN wd_in_w1[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.425 0.070 712.495 ;
    END
  END wd_in_w1[468]
  PIN wd_in_w1[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.845 0.070 712.915 ;
    END
  END wd_in_w1[469]
  PIN wd_in_w1[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 713.265 0.070 713.335 ;
    END
  END wd_in_w1[470]
  PIN wd_in_w1[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 713.685 0.070 713.755 ;
    END
  END wd_in_w1[471]
  PIN wd_in_w1[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 714.105 0.070 714.175 ;
    END
  END wd_in_w1[472]
  PIN wd_in_w1[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 714.525 0.070 714.595 ;
    END
  END wd_in_w1[473]
  PIN wd_in_w1[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 714.945 0.070 715.015 ;
    END
  END wd_in_w1[474]
  PIN wd_in_w1[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.365 0.070 715.435 ;
    END
  END wd_in_w1[475]
  PIN wd_in_w1[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.785 0.070 715.855 ;
    END
  END wd_in_w1[476]
  PIN wd_in_w1[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 716.205 0.070 716.275 ;
    END
  END wd_in_w1[477]
  PIN wd_in_w1[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 716.625 0.070 716.695 ;
    END
  END wd_in_w1[478]
  PIN wd_in_w1[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.045 0.070 717.115 ;
    END
  END wd_in_w1[479]
  PIN wd_in_w1[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.465 0.070 717.535 ;
    END
  END wd_in_w1[480]
  PIN wd_in_w1[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.885 0.070 717.955 ;
    END
  END wd_in_w1[481]
  PIN wd_in_w1[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 718.305 0.070 718.375 ;
    END
  END wd_in_w1[482]
  PIN wd_in_w1[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 718.725 0.070 718.795 ;
    END
  END wd_in_w1[483]
  PIN wd_in_w1[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.145 0.070 719.215 ;
    END
  END wd_in_w1[484]
  PIN wd_in_w1[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.565 0.070 719.635 ;
    END
  END wd_in_w1[485]
  PIN wd_in_w1[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.985 0.070 720.055 ;
    END
  END wd_in_w1[486]
  PIN wd_in_w1[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 720.405 0.070 720.475 ;
    END
  END wd_in_w1[487]
  PIN wd_in_w1[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 720.825 0.070 720.895 ;
    END
  END wd_in_w1[488]
  PIN wd_in_w1[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.245 0.070 721.315 ;
    END
  END wd_in_w1[489]
  PIN wd_in_w1[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.665 0.070 721.735 ;
    END
  END wd_in_w1[490]
  PIN wd_in_w1[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.085 0.070 722.155 ;
    END
  END wd_in_w1[491]
  PIN wd_in_w1[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.505 0.070 722.575 ;
    END
  END wd_in_w1[492]
  PIN wd_in_w1[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.925 0.070 722.995 ;
    END
  END wd_in_w1[493]
  PIN wd_in_w1[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.345 0.070 723.415 ;
    END
  END wd_in_w1[494]
  PIN wd_in_w1[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.765 0.070 723.835 ;
    END
  END wd_in_w1[495]
  PIN wd_in_w1[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.185 0.070 724.255 ;
    END
  END wd_in_w1[496]
  PIN wd_in_w1[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.605 0.070 724.675 ;
    END
  END wd_in_w1[497]
  PIN wd_in_w1[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.025 0.070 725.095 ;
    END
  END wd_in_w1[498]
  PIN wd_in_w1[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.445 0.070 725.515 ;
    END
  END wd_in_w1[499]
  PIN wd_in_w1[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.865 0.070 725.935 ;
    END
  END wd_in_w1[500]
  PIN wd_in_w1[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.285 0.070 726.355 ;
    END
  END wd_in_w1[501]
  PIN wd_in_w1[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.705 0.070 726.775 ;
    END
  END wd_in_w1[502]
  PIN wd_in_w1[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.125 0.070 727.195 ;
    END
  END wd_in_w1[503]
  PIN wd_in_w1[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.545 0.070 727.615 ;
    END
  END wd_in_w1[504]
  PIN wd_in_w1[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.965 0.070 728.035 ;
    END
  END wd_in_w1[505]
  PIN wd_in_w1[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 728.385 0.070 728.455 ;
    END
  END wd_in_w1[506]
  PIN wd_in_w1[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 728.805 0.070 728.875 ;
    END
  END wd_in_w1[507]
  PIN wd_in_w1[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.225 0.070 729.295 ;
    END
  END wd_in_w1[508]
  PIN wd_in_w1[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.645 0.070 729.715 ;
    END
  END wd_in_w1[509]
  PIN wd_in_w1[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.065 0.070 730.135 ;
    END
  END wd_in_w1[510]
  PIN wd_in_w1[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.485 0.070 730.555 ;
    END
  END wd_in_w1[511]
  PIN addr_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.045 0.070 759.115 ;
    END
  END addr_w1[0]
  PIN addr_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.465 0.070 759.535 ;
    END
  END addr_w1[1]
  PIN addr_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.885 0.070 759.955 ;
    END
  END addr_w1[2]
  PIN addr_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 760.305 0.070 760.375 ;
    END
  END addr_w1[3]
  PIN addr_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 760.725 0.070 760.795 ;
    END
  END addr_w1[4]
  PIN addr_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.145 0.070 761.215 ;
    END
  END addr_w1[5]
  PIN addr_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.565 0.070 761.635 ;
    END
  END addr_w1[6]
  PIN addr_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.985 0.070 762.055 ;
    END
  END addr_w1[7]
  PIN addr_r1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 790.545 0.070 790.615 ;
    END
  END addr_r1[0]
  PIN addr_r1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 790.965 0.070 791.035 ;
    END
  END addr_r1[1]
  PIN addr_r1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 791.385 0.070 791.455 ;
    END
  END addr_r1[2]
  PIN addr_r1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 791.805 0.070 791.875 ;
    END
  END addr_r1[3]
  PIN addr_r1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 792.225 0.070 792.295 ;
    END
  END addr_r1[4]
  PIN addr_r1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 792.645 0.070 792.715 ;
    END
  END addr_r1[5]
  PIN addr_r1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 793.065 0.070 793.135 ;
    END
  END addr_r1[6]
  PIN addr_r1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 793.485 0.070 793.555 ;
    END
  END addr_r1[7]
  PIN we_in_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 822.045 0.070 822.115 ;
    END
  END we_in_w1
  PIN ce_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 878.745 0.070 878.815 ;
    END
  END ce_w1
  PIN ce_r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 907.305 0.070 907.375 ;
    END
  END ce_r1
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 935.865 0.070 935.935 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 765.800 ;
      RECT 3.500 1.400 3.780 765.800 ;
      RECT 5.740 1.400 6.020 765.800 ;
      RECT 7.980 1.400 8.260 765.800 ;
      RECT 10.220 1.400 10.500 765.800 ;
      RECT 12.460 1.400 12.740 765.800 ;
      RECT 14.700 1.400 14.980 765.800 ;
      RECT 16.940 1.400 17.220 765.800 ;
      RECT 19.180 1.400 19.460 765.800 ;
      RECT 21.420 1.400 21.700 765.800 ;
      RECT 23.660 1.400 23.940 765.800 ;
      RECT 25.900 1.400 26.180 765.800 ;
      RECT 28.140 1.400 28.420 765.800 ;
      RECT 30.380 1.400 30.660 765.800 ;
      RECT 32.620 1.400 32.900 765.800 ;
      RECT 34.860 1.400 35.140 765.800 ;
      RECT 37.100 1.400 37.380 765.800 ;
      RECT 39.340 1.400 39.620 765.800 ;
      RECT 41.580 1.400 41.860 765.800 ;
      RECT 43.820 1.400 44.100 765.800 ;
      RECT 46.060 1.400 46.340 765.800 ;
      RECT 48.300 1.400 48.580 765.800 ;
      RECT 50.540 1.400 50.820 765.800 ;
      RECT 52.780 1.400 53.060 765.800 ;
      RECT 55.020 1.400 55.300 765.800 ;
      RECT 57.260 1.400 57.540 765.800 ;
      RECT 59.500 1.400 59.780 765.800 ;
      RECT 61.740 1.400 62.020 765.800 ;
      RECT 63.980 1.400 64.260 765.800 ;
      RECT 66.220 1.400 66.500 765.800 ;
      RECT 68.460 1.400 68.740 765.800 ;
      RECT 70.700 1.400 70.980 765.800 ;
      RECT 72.940 1.400 73.220 765.800 ;
      RECT 75.180 1.400 75.460 765.800 ;
      RECT 77.420 1.400 77.700 765.800 ;
      RECT 79.660 1.400 79.940 765.800 ;
      RECT 81.900 1.400 82.180 765.800 ;
      RECT 84.140 1.400 84.420 765.800 ;
      RECT 86.380 1.400 86.660 765.800 ;
      RECT 88.620 1.400 88.900 765.800 ;
      RECT 90.860 1.400 91.140 765.800 ;
      RECT 93.100 1.400 93.380 765.800 ;
      RECT 95.340 1.400 95.620 765.800 ;
      RECT 97.580 1.400 97.860 765.800 ;
      RECT 99.820 1.400 100.100 765.800 ;
      RECT 102.060 1.400 102.340 765.800 ;
      RECT 104.300 1.400 104.580 765.800 ;
      RECT 106.540 1.400 106.820 765.800 ;
      RECT 108.780 1.400 109.060 765.800 ;
      RECT 111.020 1.400 111.300 765.800 ;
      RECT 113.260 1.400 113.540 765.800 ;
      RECT 115.500 1.400 115.780 765.800 ;
      RECT 117.740 1.400 118.020 765.800 ;
      RECT 119.980 1.400 120.260 765.800 ;
      RECT 122.220 1.400 122.500 765.800 ;
      RECT 124.460 1.400 124.740 765.800 ;
      RECT 126.700 1.400 126.980 765.800 ;
      RECT 128.940 1.400 129.220 765.800 ;
      RECT 131.180 1.400 131.460 765.800 ;
      RECT 133.420 1.400 133.700 765.800 ;
      RECT 135.660 1.400 135.940 765.800 ;
      RECT 137.900 1.400 138.180 765.800 ;
      RECT 140.140 1.400 140.420 765.800 ;
      RECT 142.380 1.400 142.660 765.800 ;
      RECT 144.620 1.400 144.900 765.800 ;
      RECT 146.860 1.400 147.140 765.800 ;
      RECT 149.100 1.400 149.380 765.800 ;
      RECT 151.340 1.400 151.620 765.800 ;
      RECT 153.580 1.400 153.860 765.800 ;
      RECT 155.820 1.400 156.100 765.800 ;
      RECT 158.060 1.400 158.340 765.800 ;
      RECT 160.300 1.400 160.580 765.800 ;
      RECT 162.540 1.400 162.820 765.800 ;
      RECT 164.780 1.400 165.060 765.800 ;
      RECT 167.020 1.400 167.300 765.800 ;
      RECT 169.260 1.400 169.540 765.800 ;
      RECT 171.500 1.400 171.780 765.800 ;
      RECT 173.740 1.400 174.020 765.800 ;
      RECT 175.980 1.400 176.260 765.800 ;
      RECT 178.220 1.400 178.500 765.800 ;
      RECT 180.460 1.400 180.740 765.800 ;
      RECT 182.700 1.400 182.980 765.800 ;
      RECT 184.940 1.400 185.220 765.800 ;
      RECT 187.180 1.400 187.460 765.800 ;
      RECT 189.420 1.400 189.700 765.800 ;
      RECT 191.660 1.400 191.940 765.800 ;
      RECT 193.900 1.400 194.180 765.800 ;
      RECT 196.140 1.400 196.420 765.800 ;
      RECT 198.380 1.400 198.660 765.800 ;
      RECT 200.620 1.400 200.900 765.800 ;
      RECT 202.860 1.400 203.140 765.800 ;
      RECT 205.100 1.400 205.380 765.800 ;
      RECT 207.340 1.400 207.620 765.800 ;
      RECT 209.580 1.400 209.860 765.800 ;
      RECT 211.820 1.400 212.100 765.800 ;
      RECT 214.060 1.400 214.340 765.800 ;
      RECT 216.300 1.400 216.580 765.800 ;
      RECT 218.540 1.400 218.820 765.800 ;
      RECT 220.780 1.400 221.060 765.800 ;
      RECT 223.020 1.400 223.300 765.800 ;
      RECT 225.260 1.400 225.540 765.800 ;
      RECT 227.500 1.400 227.780 765.800 ;
      RECT 229.740 1.400 230.020 765.800 ;
      RECT 231.980 1.400 232.260 765.800 ;
      RECT 234.220 1.400 234.500 765.800 ;
      RECT 236.460 1.400 236.740 765.800 ;
      RECT 238.700 1.400 238.980 765.800 ;
      RECT 240.940 1.400 241.220 765.800 ;
      RECT 243.180 1.400 243.460 765.800 ;
      RECT 245.420 1.400 245.700 765.800 ;
      RECT 247.660 1.400 247.940 765.800 ;
      RECT 249.900 1.400 250.180 765.800 ;
      RECT 252.140 1.400 252.420 765.800 ;
      RECT 254.380 1.400 254.660 765.800 ;
      RECT 256.620 1.400 256.900 765.800 ;
      RECT 258.860 1.400 259.140 765.800 ;
      RECT 261.100 1.400 261.380 765.800 ;
      RECT 263.340 1.400 263.620 765.800 ;
      RECT 265.580 1.400 265.860 765.800 ;
      RECT 267.820 1.400 268.100 765.800 ;
      RECT 270.060 1.400 270.340 765.800 ;
      RECT 272.300 1.400 272.580 765.800 ;
      RECT 274.540 1.400 274.820 765.800 ;
      RECT 276.780 1.400 277.060 765.800 ;
      RECT 279.020 1.400 279.300 765.800 ;
      RECT 281.260 1.400 281.540 765.800 ;
      RECT 283.500 1.400 283.780 765.800 ;
      RECT 285.740 1.400 286.020 765.800 ;
      RECT 287.980 1.400 288.260 765.800 ;
      RECT 290.220 1.400 290.500 765.800 ;
      RECT 292.460 1.400 292.740 765.800 ;
      RECT 294.700 1.400 294.980 765.800 ;
      RECT 296.940 1.400 297.220 765.800 ;
      RECT 299.180 1.400 299.460 765.800 ;
      RECT 301.420 1.400 301.700 765.800 ;
      RECT 303.660 1.400 303.940 765.800 ;
      RECT 305.900 1.400 306.180 765.800 ;
      RECT 308.140 1.400 308.420 765.800 ;
      RECT 310.380 1.400 310.660 765.800 ;
      RECT 312.620 1.400 312.900 765.800 ;
      RECT 314.860 1.400 315.140 765.800 ;
      RECT 317.100 1.400 317.380 765.800 ;
      RECT 319.340 1.400 319.620 765.800 ;
      RECT 321.580 1.400 321.860 765.800 ;
      RECT 323.820 1.400 324.100 765.800 ;
      RECT 326.060 1.400 326.340 765.800 ;
      RECT 328.300 1.400 328.580 765.800 ;
      RECT 330.540 1.400 330.820 765.800 ;
      RECT 332.780 1.400 333.060 765.800 ;
      RECT 335.020 1.400 335.300 765.800 ;
      RECT 337.260 1.400 337.540 765.800 ;
      RECT 339.500 1.400 339.780 765.800 ;
      RECT 341.740 1.400 342.020 765.800 ;
      RECT 343.980 1.400 344.260 765.800 ;
      RECT 346.220 1.400 346.500 765.800 ;
      RECT 348.460 1.400 348.740 765.800 ;
      RECT 350.700 1.400 350.980 765.800 ;
      RECT 352.940 1.400 353.220 765.800 ;
      RECT 355.180 1.400 355.460 765.800 ;
      RECT 357.420 1.400 357.700 765.800 ;
      RECT 359.660 1.400 359.940 765.800 ;
      RECT 361.900 1.400 362.180 765.800 ;
      RECT 364.140 1.400 364.420 765.800 ;
      RECT 366.380 1.400 366.660 765.800 ;
      RECT 368.620 1.400 368.900 765.800 ;
      RECT 370.860 1.400 371.140 765.800 ;
      RECT 373.100 1.400 373.380 765.800 ;
      RECT 375.340 1.400 375.620 765.800 ;
      RECT 377.580 1.400 377.860 765.800 ;
      RECT 379.820 1.400 380.100 765.800 ;
      RECT 382.060 1.400 382.340 765.800 ;
      RECT 384.300 1.400 384.580 765.800 ;
      RECT 386.540 1.400 386.820 765.800 ;
      RECT 388.780 1.400 389.060 765.800 ;
      RECT 391.020 1.400 391.300 765.800 ;
      RECT 393.260 1.400 393.540 765.800 ;
      RECT 395.500 1.400 395.780 765.800 ;
      RECT 397.740 1.400 398.020 765.800 ;
      RECT 399.980 1.400 400.260 765.800 ;
      RECT 402.220 1.400 402.500 765.800 ;
      RECT 404.460 1.400 404.740 765.800 ;
      RECT 406.700 1.400 406.980 765.800 ;
      RECT 408.940 1.400 409.220 765.800 ;
      RECT 411.180 1.400 411.460 765.800 ;
      RECT 413.420 1.400 413.700 765.800 ;
      RECT 415.660 1.400 415.940 765.800 ;
      RECT 417.900 1.400 418.180 765.800 ;
      RECT 420.140 1.400 420.420 765.800 ;
      RECT 422.380 1.400 422.660 765.800 ;
      RECT 424.620 1.400 424.900 765.800 ;
      RECT 426.860 1.400 427.140 765.800 ;
      RECT 429.100 1.400 429.380 765.800 ;
      RECT 431.340 1.400 431.620 765.800 ;
      RECT 433.580 1.400 433.860 765.800 ;
      RECT 435.820 1.400 436.100 765.800 ;
      RECT 438.060 1.400 438.340 765.800 ;
      RECT 440.300 1.400 440.580 765.800 ;
      RECT 442.540 1.400 442.820 765.800 ;
      RECT 444.780 1.400 445.060 765.800 ;
      RECT 447.020 1.400 447.300 765.800 ;
      RECT 449.260 1.400 449.540 765.800 ;
      RECT 451.500 1.400 451.780 765.800 ;
      RECT 453.740 1.400 454.020 765.800 ;
      RECT 455.980 1.400 456.260 765.800 ;
      RECT 458.220 1.400 458.500 765.800 ;
      RECT 460.460 1.400 460.740 765.800 ;
      RECT 462.700 1.400 462.980 765.800 ;
      RECT 464.940 1.400 465.220 765.800 ;
      RECT 467.180 1.400 467.460 765.800 ;
      RECT 469.420 1.400 469.700 765.800 ;
      RECT 471.660 1.400 471.940 765.800 ;
      RECT 473.900 1.400 474.180 765.800 ;
      RECT 476.140 1.400 476.420 765.800 ;
      RECT 478.380 1.400 478.660 765.800 ;
      RECT 480.620 1.400 480.900 765.800 ;
      RECT 482.860 1.400 483.140 765.800 ;
      RECT 485.100 1.400 485.380 765.800 ;
      RECT 487.340 1.400 487.620 765.800 ;
      RECT 489.580 1.400 489.860 765.800 ;
      RECT 491.820 1.400 492.100 765.800 ;
      RECT 494.060 1.400 494.340 765.800 ;
      RECT 496.300 1.400 496.580 765.800 ;
      RECT 498.540 1.400 498.820 765.800 ;
      RECT 500.780 1.400 501.060 765.800 ;
      RECT 503.020 1.400 503.300 765.800 ;
      RECT 505.260 1.400 505.540 765.800 ;
      RECT 507.500 1.400 507.780 765.800 ;
      RECT 509.740 1.400 510.020 765.800 ;
      RECT 511.980 1.400 512.260 765.800 ;
      RECT 514.220 1.400 514.500 765.800 ;
      RECT 516.460 1.400 516.740 765.800 ;
      RECT 518.700 1.400 518.980 765.800 ;
      RECT 520.940 1.400 521.220 765.800 ;
      RECT 523.180 1.400 523.460 765.800 ;
      RECT 525.420 1.400 525.700 765.800 ;
      RECT 527.660 1.400 527.940 765.800 ;
      RECT 529.900 1.400 530.180 765.800 ;
      RECT 532.140 1.400 532.420 765.800 ;
      RECT 534.380 1.400 534.660 765.800 ;
      RECT 536.620 1.400 536.900 765.800 ;
      RECT 538.860 1.400 539.140 765.800 ;
      RECT 541.100 1.400 541.380 765.800 ;
      RECT 543.340 1.400 543.620 765.800 ;
      RECT 545.580 1.400 545.860 765.800 ;
      RECT 547.820 1.400 548.100 765.800 ;
      RECT 550.060 1.400 550.340 765.800 ;
      RECT 552.300 1.400 552.580 765.800 ;
      RECT 554.540 1.400 554.820 765.800 ;
      RECT 556.780 1.400 557.060 765.800 ;
      RECT 559.020 1.400 559.300 765.800 ;
      RECT 561.260 1.400 561.540 765.800 ;
      RECT 563.500 1.400 563.780 765.800 ;
      RECT 565.740 1.400 566.020 765.800 ;
      RECT 567.980 1.400 568.260 765.800 ;
      RECT 570.220 1.400 570.500 765.800 ;
      RECT 572.460 1.400 572.740 765.800 ;
      RECT 574.700 1.400 574.980 765.800 ;
      RECT 576.940 1.400 577.220 765.800 ;
      RECT 579.180 1.400 579.460 765.800 ;
      RECT 581.420 1.400 581.700 765.800 ;
      RECT 583.660 1.400 583.940 765.800 ;
      RECT 585.900 1.400 586.180 765.800 ;
      RECT 588.140 1.400 588.420 765.800 ;
      RECT 590.380 1.400 590.660 765.800 ;
      RECT 592.620 1.400 592.900 765.800 ;
      RECT 594.860 1.400 595.140 765.800 ;
      RECT 597.100 1.400 597.380 765.800 ;
      RECT 599.340 1.400 599.620 765.800 ;
      RECT 601.580 1.400 601.860 765.800 ;
      RECT 603.820 1.400 604.100 765.800 ;
      RECT 606.060 1.400 606.340 765.800 ;
      RECT 608.300 1.400 608.580 765.800 ;
      RECT 610.540 1.400 610.820 765.800 ;
      RECT 612.780 1.400 613.060 765.800 ;
      RECT 615.020 1.400 615.300 765.800 ;
      RECT 617.260 1.400 617.540 765.800 ;
      RECT 619.500 1.400 619.780 765.800 ;
      RECT 621.740 1.400 622.020 765.800 ;
      RECT 623.980 1.400 624.260 765.800 ;
      RECT 626.220 1.400 626.500 765.800 ;
      RECT 628.460 1.400 628.740 765.800 ;
      RECT 630.700 1.400 630.980 765.800 ;
      RECT 632.940 1.400 633.220 765.800 ;
      RECT 635.180 1.400 635.460 765.800 ;
      RECT 637.420 1.400 637.700 765.800 ;
      RECT 639.660 1.400 639.940 765.800 ;
      RECT 641.900 1.400 642.180 765.800 ;
      RECT 644.140 1.400 644.420 765.800 ;
      RECT 646.380 1.400 646.660 765.800 ;
      RECT 648.620 1.400 648.900 765.800 ;
      RECT 650.860 1.400 651.140 765.800 ;
      RECT 653.100 1.400 653.380 765.800 ;
      RECT 655.340 1.400 655.620 765.800 ;
      RECT 657.580 1.400 657.860 765.800 ;
      RECT 659.820 1.400 660.100 765.800 ;
      RECT 662.060 1.400 662.340 765.800 ;
      RECT 664.300 1.400 664.580 765.800 ;
      RECT 666.540 1.400 666.820 765.800 ;
      RECT 668.780 1.400 669.060 765.800 ;
      RECT 671.020 1.400 671.300 765.800 ;
      RECT 673.260 1.400 673.540 765.800 ;
      RECT 675.500 1.400 675.780 765.800 ;
      RECT 677.740 1.400 678.020 765.800 ;
      RECT 679.980 1.400 680.260 765.800 ;
      RECT 682.220 1.400 682.500 765.800 ;
      RECT 684.460 1.400 684.740 765.800 ;
      RECT 686.700 1.400 686.980 765.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 765.800 ;
      RECT 4.620 1.400 4.900 765.800 ;
      RECT 6.860 1.400 7.140 765.800 ;
      RECT 9.100 1.400 9.380 765.800 ;
      RECT 11.340 1.400 11.620 765.800 ;
      RECT 13.580 1.400 13.860 765.800 ;
      RECT 15.820 1.400 16.100 765.800 ;
      RECT 18.060 1.400 18.340 765.800 ;
      RECT 20.300 1.400 20.580 765.800 ;
      RECT 22.540 1.400 22.820 765.800 ;
      RECT 24.780 1.400 25.060 765.800 ;
      RECT 27.020 1.400 27.300 765.800 ;
      RECT 29.260 1.400 29.540 765.800 ;
      RECT 31.500 1.400 31.780 765.800 ;
      RECT 33.740 1.400 34.020 765.800 ;
      RECT 35.980 1.400 36.260 765.800 ;
      RECT 38.220 1.400 38.500 765.800 ;
      RECT 40.460 1.400 40.740 765.800 ;
      RECT 42.700 1.400 42.980 765.800 ;
      RECT 44.940 1.400 45.220 765.800 ;
      RECT 47.180 1.400 47.460 765.800 ;
      RECT 49.420 1.400 49.700 765.800 ;
      RECT 51.660 1.400 51.940 765.800 ;
      RECT 53.900 1.400 54.180 765.800 ;
      RECT 56.140 1.400 56.420 765.800 ;
      RECT 58.380 1.400 58.660 765.800 ;
      RECT 60.620 1.400 60.900 765.800 ;
      RECT 62.860 1.400 63.140 765.800 ;
      RECT 65.100 1.400 65.380 765.800 ;
      RECT 67.340 1.400 67.620 765.800 ;
      RECT 69.580 1.400 69.860 765.800 ;
      RECT 71.820 1.400 72.100 765.800 ;
      RECT 74.060 1.400 74.340 765.800 ;
      RECT 76.300 1.400 76.580 765.800 ;
      RECT 78.540 1.400 78.820 765.800 ;
      RECT 80.780 1.400 81.060 765.800 ;
      RECT 83.020 1.400 83.300 765.800 ;
      RECT 85.260 1.400 85.540 765.800 ;
      RECT 87.500 1.400 87.780 765.800 ;
      RECT 89.740 1.400 90.020 765.800 ;
      RECT 91.980 1.400 92.260 765.800 ;
      RECT 94.220 1.400 94.500 765.800 ;
      RECT 96.460 1.400 96.740 765.800 ;
      RECT 98.700 1.400 98.980 765.800 ;
      RECT 100.940 1.400 101.220 765.800 ;
      RECT 103.180 1.400 103.460 765.800 ;
      RECT 105.420 1.400 105.700 765.800 ;
      RECT 107.660 1.400 107.940 765.800 ;
      RECT 109.900 1.400 110.180 765.800 ;
      RECT 112.140 1.400 112.420 765.800 ;
      RECT 114.380 1.400 114.660 765.800 ;
      RECT 116.620 1.400 116.900 765.800 ;
      RECT 118.860 1.400 119.140 765.800 ;
      RECT 121.100 1.400 121.380 765.800 ;
      RECT 123.340 1.400 123.620 765.800 ;
      RECT 125.580 1.400 125.860 765.800 ;
      RECT 127.820 1.400 128.100 765.800 ;
      RECT 130.060 1.400 130.340 765.800 ;
      RECT 132.300 1.400 132.580 765.800 ;
      RECT 134.540 1.400 134.820 765.800 ;
      RECT 136.780 1.400 137.060 765.800 ;
      RECT 139.020 1.400 139.300 765.800 ;
      RECT 141.260 1.400 141.540 765.800 ;
      RECT 143.500 1.400 143.780 765.800 ;
      RECT 145.740 1.400 146.020 765.800 ;
      RECT 147.980 1.400 148.260 765.800 ;
      RECT 150.220 1.400 150.500 765.800 ;
      RECT 152.460 1.400 152.740 765.800 ;
      RECT 154.700 1.400 154.980 765.800 ;
      RECT 156.940 1.400 157.220 765.800 ;
      RECT 159.180 1.400 159.460 765.800 ;
      RECT 161.420 1.400 161.700 765.800 ;
      RECT 163.660 1.400 163.940 765.800 ;
      RECT 165.900 1.400 166.180 765.800 ;
      RECT 168.140 1.400 168.420 765.800 ;
      RECT 170.380 1.400 170.660 765.800 ;
      RECT 172.620 1.400 172.900 765.800 ;
      RECT 174.860 1.400 175.140 765.800 ;
      RECT 177.100 1.400 177.380 765.800 ;
      RECT 179.340 1.400 179.620 765.800 ;
      RECT 181.580 1.400 181.860 765.800 ;
      RECT 183.820 1.400 184.100 765.800 ;
      RECT 186.060 1.400 186.340 765.800 ;
      RECT 188.300 1.400 188.580 765.800 ;
      RECT 190.540 1.400 190.820 765.800 ;
      RECT 192.780 1.400 193.060 765.800 ;
      RECT 195.020 1.400 195.300 765.800 ;
      RECT 197.260 1.400 197.540 765.800 ;
      RECT 199.500 1.400 199.780 765.800 ;
      RECT 201.740 1.400 202.020 765.800 ;
      RECT 203.980 1.400 204.260 765.800 ;
      RECT 206.220 1.400 206.500 765.800 ;
      RECT 208.460 1.400 208.740 765.800 ;
      RECT 210.700 1.400 210.980 765.800 ;
      RECT 212.940 1.400 213.220 765.800 ;
      RECT 215.180 1.400 215.460 765.800 ;
      RECT 217.420 1.400 217.700 765.800 ;
      RECT 219.660 1.400 219.940 765.800 ;
      RECT 221.900 1.400 222.180 765.800 ;
      RECT 224.140 1.400 224.420 765.800 ;
      RECT 226.380 1.400 226.660 765.800 ;
      RECT 228.620 1.400 228.900 765.800 ;
      RECT 230.860 1.400 231.140 765.800 ;
      RECT 233.100 1.400 233.380 765.800 ;
      RECT 235.340 1.400 235.620 765.800 ;
      RECT 237.580 1.400 237.860 765.800 ;
      RECT 239.820 1.400 240.100 765.800 ;
      RECT 242.060 1.400 242.340 765.800 ;
      RECT 244.300 1.400 244.580 765.800 ;
      RECT 246.540 1.400 246.820 765.800 ;
      RECT 248.780 1.400 249.060 765.800 ;
      RECT 251.020 1.400 251.300 765.800 ;
      RECT 253.260 1.400 253.540 765.800 ;
      RECT 255.500 1.400 255.780 765.800 ;
      RECT 257.740 1.400 258.020 765.800 ;
      RECT 259.980 1.400 260.260 765.800 ;
      RECT 262.220 1.400 262.500 765.800 ;
      RECT 264.460 1.400 264.740 765.800 ;
      RECT 266.700 1.400 266.980 765.800 ;
      RECT 268.940 1.400 269.220 765.800 ;
      RECT 271.180 1.400 271.460 765.800 ;
      RECT 273.420 1.400 273.700 765.800 ;
      RECT 275.660 1.400 275.940 765.800 ;
      RECT 277.900 1.400 278.180 765.800 ;
      RECT 280.140 1.400 280.420 765.800 ;
      RECT 282.380 1.400 282.660 765.800 ;
      RECT 284.620 1.400 284.900 765.800 ;
      RECT 286.860 1.400 287.140 765.800 ;
      RECT 289.100 1.400 289.380 765.800 ;
      RECT 291.340 1.400 291.620 765.800 ;
      RECT 293.580 1.400 293.860 765.800 ;
      RECT 295.820 1.400 296.100 765.800 ;
      RECT 298.060 1.400 298.340 765.800 ;
      RECT 300.300 1.400 300.580 765.800 ;
      RECT 302.540 1.400 302.820 765.800 ;
      RECT 304.780 1.400 305.060 765.800 ;
      RECT 307.020 1.400 307.300 765.800 ;
      RECT 309.260 1.400 309.540 765.800 ;
      RECT 311.500 1.400 311.780 765.800 ;
      RECT 313.740 1.400 314.020 765.800 ;
      RECT 315.980 1.400 316.260 765.800 ;
      RECT 318.220 1.400 318.500 765.800 ;
      RECT 320.460 1.400 320.740 765.800 ;
      RECT 322.700 1.400 322.980 765.800 ;
      RECT 324.940 1.400 325.220 765.800 ;
      RECT 327.180 1.400 327.460 765.800 ;
      RECT 329.420 1.400 329.700 765.800 ;
      RECT 331.660 1.400 331.940 765.800 ;
      RECT 333.900 1.400 334.180 765.800 ;
      RECT 336.140 1.400 336.420 765.800 ;
      RECT 338.380 1.400 338.660 765.800 ;
      RECT 340.620 1.400 340.900 765.800 ;
      RECT 342.860 1.400 343.140 765.800 ;
      RECT 345.100 1.400 345.380 765.800 ;
      RECT 347.340 1.400 347.620 765.800 ;
      RECT 349.580 1.400 349.860 765.800 ;
      RECT 351.820 1.400 352.100 765.800 ;
      RECT 354.060 1.400 354.340 765.800 ;
      RECT 356.300 1.400 356.580 765.800 ;
      RECT 358.540 1.400 358.820 765.800 ;
      RECT 360.780 1.400 361.060 765.800 ;
      RECT 363.020 1.400 363.300 765.800 ;
      RECT 365.260 1.400 365.540 765.800 ;
      RECT 367.500 1.400 367.780 765.800 ;
      RECT 369.740 1.400 370.020 765.800 ;
      RECT 371.980 1.400 372.260 765.800 ;
      RECT 374.220 1.400 374.500 765.800 ;
      RECT 376.460 1.400 376.740 765.800 ;
      RECT 378.700 1.400 378.980 765.800 ;
      RECT 380.940 1.400 381.220 765.800 ;
      RECT 383.180 1.400 383.460 765.800 ;
      RECT 385.420 1.400 385.700 765.800 ;
      RECT 387.660 1.400 387.940 765.800 ;
      RECT 389.900 1.400 390.180 765.800 ;
      RECT 392.140 1.400 392.420 765.800 ;
      RECT 394.380 1.400 394.660 765.800 ;
      RECT 396.620 1.400 396.900 765.800 ;
      RECT 398.860 1.400 399.140 765.800 ;
      RECT 401.100 1.400 401.380 765.800 ;
      RECT 403.340 1.400 403.620 765.800 ;
      RECT 405.580 1.400 405.860 765.800 ;
      RECT 407.820 1.400 408.100 765.800 ;
      RECT 410.060 1.400 410.340 765.800 ;
      RECT 412.300 1.400 412.580 765.800 ;
      RECT 414.540 1.400 414.820 765.800 ;
      RECT 416.780 1.400 417.060 765.800 ;
      RECT 419.020 1.400 419.300 765.800 ;
      RECT 421.260 1.400 421.540 765.800 ;
      RECT 423.500 1.400 423.780 765.800 ;
      RECT 425.740 1.400 426.020 765.800 ;
      RECT 427.980 1.400 428.260 765.800 ;
      RECT 430.220 1.400 430.500 765.800 ;
      RECT 432.460 1.400 432.740 765.800 ;
      RECT 434.700 1.400 434.980 765.800 ;
      RECT 436.940 1.400 437.220 765.800 ;
      RECT 439.180 1.400 439.460 765.800 ;
      RECT 441.420 1.400 441.700 765.800 ;
      RECT 443.660 1.400 443.940 765.800 ;
      RECT 445.900 1.400 446.180 765.800 ;
      RECT 448.140 1.400 448.420 765.800 ;
      RECT 450.380 1.400 450.660 765.800 ;
      RECT 452.620 1.400 452.900 765.800 ;
      RECT 454.860 1.400 455.140 765.800 ;
      RECT 457.100 1.400 457.380 765.800 ;
      RECT 459.340 1.400 459.620 765.800 ;
      RECT 461.580 1.400 461.860 765.800 ;
      RECT 463.820 1.400 464.100 765.800 ;
      RECT 466.060 1.400 466.340 765.800 ;
      RECT 468.300 1.400 468.580 765.800 ;
      RECT 470.540 1.400 470.820 765.800 ;
      RECT 472.780 1.400 473.060 765.800 ;
      RECT 475.020 1.400 475.300 765.800 ;
      RECT 477.260 1.400 477.540 765.800 ;
      RECT 479.500 1.400 479.780 765.800 ;
      RECT 481.740 1.400 482.020 765.800 ;
      RECT 483.980 1.400 484.260 765.800 ;
      RECT 486.220 1.400 486.500 765.800 ;
      RECT 488.460 1.400 488.740 765.800 ;
      RECT 490.700 1.400 490.980 765.800 ;
      RECT 492.940 1.400 493.220 765.800 ;
      RECT 495.180 1.400 495.460 765.800 ;
      RECT 497.420 1.400 497.700 765.800 ;
      RECT 499.660 1.400 499.940 765.800 ;
      RECT 501.900 1.400 502.180 765.800 ;
      RECT 504.140 1.400 504.420 765.800 ;
      RECT 506.380 1.400 506.660 765.800 ;
      RECT 508.620 1.400 508.900 765.800 ;
      RECT 510.860 1.400 511.140 765.800 ;
      RECT 513.100 1.400 513.380 765.800 ;
      RECT 515.340 1.400 515.620 765.800 ;
      RECT 517.580 1.400 517.860 765.800 ;
      RECT 519.820 1.400 520.100 765.800 ;
      RECT 522.060 1.400 522.340 765.800 ;
      RECT 524.300 1.400 524.580 765.800 ;
      RECT 526.540 1.400 526.820 765.800 ;
      RECT 528.780 1.400 529.060 765.800 ;
      RECT 531.020 1.400 531.300 765.800 ;
      RECT 533.260 1.400 533.540 765.800 ;
      RECT 535.500 1.400 535.780 765.800 ;
      RECT 537.740 1.400 538.020 765.800 ;
      RECT 539.980 1.400 540.260 765.800 ;
      RECT 542.220 1.400 542.500 765.800 ;
      RECT 544.460 1.400 544.740 765.800 ;
      RECT 546.700 1.400 546.980 765.800 ;
      RECT 548.940 1.400 549.220 765.800 ;
      RECT 551.180 1.400 551.460 765.800 ;
      RECT 553.420 1.400 553.700 765.800 ;
      RECT 555.660 1.400 555.940 765.800 ;
      RECT 557.900 1.400 558.180 765.800 ;
      RECT 560.140 1.400 560.420 765.800 ;
      RECT 562.380 1.400 562.660 765.800 ;
      RECT 564.620 1.400 564.900 765.800 ;
      RECT 566.860 1.400 567.140 765.800 ;
      RECT 569.100 1.400 569.380 765.800 ;
      RECT 571.340 1.400 571.620 765.800 ;
      RECT 573.580 1.400 573.860 765.800 ;
      RECT 575.820 1.400 576.100 765.800 ;
      RECT 578.060 1.400 578.340 765.800 ;
      RECT 580.300 1.400 580.580 765.800 ;
      RECT 582.540 1.400 582.820 765.800 ;
      RECT 584.780 1.400 585.060 765.800 ;
      RECT 587.020 1.400 587.300 765.800 ;
      RECT 589.260 1.400 589.540 765.800 ;
      RECT 591.500 1.400 591.780 765.800 ;
      RECT 593.740 1.400 594.020 765.800 ;
      RECT 595.980 1.400 596.260 765.800 ;
      RECT 598.220 1.400 598.500 765.800 ;
      RECT 600.460 1.400 600.740 765.800 ;
      RECT 602.700 1.400 602.980 765.800 ;
      RECT 604.940 1.400 605.220 765.800 ;
      RECT 607.180 1.400 607.460 765.800 ;
      RECT 609.420 1.400 609.700 765.800 ;
      RECT 611.660 1.400 611.940 765.800 ;
      RECT 613.900 1.400 614.180 765.800 ;
      RECT 616.140 1.400 616.420 765.800 ;
      RECT 618.380 1.400 618.660 765.800 ;
      RECT 620.620 1.400 620.900 765.800 ;
      RECT 622.860 1.400 623.140 765.800 ;
      RECT 625.100 1.400 625.380 765.800 ;
      RECT 627.340 1.400 627.620 765.800 ;
      RECT 629.580 1.400 629.860 765.800 ;
      RECT 631.820 1.400 632.100 765.800 ;
      RECT 634.060 1.400 634.340 765.800 ;
      RECT 636.300 1.400 636.580 765.800 ;
      RECT 638.540 1.400 638.820 765.800 ;
      RECT 640.780 1.400 641.060 765.800 ;
      RECT 643.020 1.400 643.300 765.800 ;
      RECT 645.260 1.400 645.540 765.800 ;
      RECT 647.500 1.400 647.780 765.800 ;
      RECT 649.740 1.400 650.020 765.800 ;
      RECT 651.980 1.400 652.260 765.800 ;
      RECT 654.220 1.400 654.500 765.800 ;
      RECT 656.460 1.400 656.740 765.800 ;
      RECT 658.700 1.400 658.980 765.800 ;
      RECT 660.940 1.400 661.220 765.800 ;
      RECT 663.180 1.400 663.460 765.800 ;
      RECT 665.420 1.400 665.700 765.800 ;
      RECT 667.660 1.400 667.940 765.800 ;
      RECT 669.900 1.400 670.180 765.800 ;
      RECT 672.140 1.400 672.420 765.800 ;
      RECT 674.380 1.400 674.660 765.800 ;
      RECT 676.620 1.400 676.900 765.800 ;
      RECT 678.860 1.400 679.140 765.800 ;
      RECT 681.100 1.400 681.380 765.800 ;
      RECT 683.340 1.400 683.620 765.800 ;
      RECT 685.580 1.400 685.860 765.800 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 689.130 767.200 ;
    LAYER metal2 ;
    RECT 0 0 689.130 767.200 ;
    LAYER metal3 ;
    RECT 0.070 0 689.130 767.200 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.785 ;
    RECT 0 1.855 0.070 2.205 ;
    RECT 0 2.275 0.070 2.625 ;
    RECT 0 2.695 0.070 3.045 ;
    RECT 0 3.115 0.070 3.465 ;
    RECT 0 3.535 0.070 3.885 ;
    RECT 0 3.955 0.070 4.305 ;
    RECT 0 4.375 0.070 4.725 ;
    RECT 0 4.795 0.070 5.145 ;
    RECT 0 5.215 0.070 5.565 ;
    RECT 0 5.635 0.070 5.985 ;
    RECT 0 6.055 0.070 6.405 ;
    RECT 0 6.475 0.070 6.825 ;
    RECT 0 6.895 0.070 7.245 ;
    RECT 0 7.315 0.070 7.665 ;
    RECT 0 7.735 0.070 8.085 ;
    RECT 0 8.155 0.070 8.505 ;
    RECT 0 8.575 0.070 8.925 ;
    RECT 0 8.995 0.070 9.345 ;
    RECT 0 9.415 0.070 9.765 ;
    RECT 0 9.835 0.070 10.185 ;
    RECT 0 10.255 0.070 10.605 ;
    RECT 0 10.675 0.070 11.025 ;
    RECT 0 11.095 0.070 11.445 ;
    RECT 0 11.515 0.070 11.865 ;
    RECT 0 11.935 0.070 12.285 ;
    RECT 0 12.355 0.070 12.705 ;
    RECT 0 12.775 0.070 13.125 ;
    RECT 0 13.195 0.070 13.545 ;
    RECT 0 13.615 0.070 13.965 ;
    RECT 0 14.035 0.070 14.385 ;
    RECT 0 14.455 0.070 14.805 ;
    RECT 0 14.875 0.070 15.225 ;
    RECT 0 15.295 0.070 15.645 ;
    RECT 0 15.715 0.070 16.065 ;
    RECT 0 16.135 0.070 16.485 ;
    RECT 0 16.555 0.070 16.905 ;
    RECT 0 16.975 0.070 17.325 ;
    RECT 0 17.395 0.070 17.745 ;
    RECT 0 17.815 0.070 18.165 ;
    RECT 0 18.235 0.070 18.585 ;
    RECT 0 18.655 0.070 19.005 ;
    RECT 0 19.075 0.070 19.425 ;
    RECT 0 19.495 0.070 19.845 ;
    RECT 0 19.915 0.070 20.265 ;
    RECT 0 20.335 0.070 20.685 ;
    RECT 0 20.755 0.070 21.105 ;
    RECT 0 21.175 0.070 21.525 ;
    RECT 0 21.595 0.070 21.945 ;
    RECT 0 22.015 0.070 22.365 ;
    RECT 0 22.435 0.070 22.785 ;
    RECT 0 22.855 0.070 23.205 ;
    RECT 0 23.275 0.070 23.625 ;
    RECT 0 23.695 0.070 24.045 ;
    RECT 0 24.115 0.070 24.465 ;
    RECT 0 24.535 0.070 24.885 ;
    RECT 0 24.955 0.070 25.305 ;
    RECT 0 25.375 0.070 25.725 ;
    RECT 0 25.795 0.070 26.145 ;
    RECT 0 26.215 0.070 26.565 ;
    RECT 0 26.635 0.070 26.985 ;
    RECT 0 27.055 0.070 27.405 ;
    RECT 0 27.475 0.070 27.825 ;
    RECT 0 27.895 0.070 28.245 ;
    RECT 0 28.315 0.070 28.665 ;
    RECT 0 28.735 0.070 29.085 ;
    RECT 0 29.155 0.070 29.505 ;
    RECT 0 29.575 0.070 29.925 ;
    RECT 0 29.995 0.070 30.345 ;
    RECT 0 30.415 0.070 30.765 ;
    RECT 0 30.835 0.070 31.185 ;
    RECT 0 31.255 0.070 31.605 ;
    RECT 0 31.675 0.070 32.025 ;
    RECT 0 32.095 0.070 32.445 ;
    RECT 0 32.515 0.070 32.865 ;
    RECT 0 32.935 0.070 33.285 ;
    RECT 0 33.355 0.070 33.705 ;
    RECT 0 33.775 0.070 34.125 ;
    RECT 0 34.195 0.070 34.545 ;
    RECT 0 34.615 0.070 34.965 ;
    RECT 0 35.035 0.070 35.385 ;
    RECT 0 35.455 0.070 35.805 ;
    RECT 0 35.875 0.070 36.225 ;
    RECT 0 36.295 0.070 36.645 ;
    RECT 0 36.715 0.070 37.065 ;
    RECT 0 37.135 0.070 37.485 ;
    RECT 0 37.555 0.070 37.905 ;
    RECT 0 37.975 0.070 38.325 ;
    RECT 0 38.395 0.070 38.745 ;
    RECT 0 38.815 0.070 39.165 ;
    RECT 0 39.235 0.070 39.585 ;
    RECT 0 39.655 0.070 40.005 ;
    RECT 0 40.075 0.070 40.425 ;
    RECT 0 40.495 0.070 40.845 ;
    RECT 0 40.915 0.070 41.265 ;
    RECT 0 41.335 0.070 41.685 ;
    RECT 0 41.755 0.070 42.105 ;
    RECT 0 42.175 0.070 42.525 ;
    RECT 0 42.595 0.070 42.945 ;
    RECT 0 43.015 0.070 43.365 ;
    RECT 0 43.435 0.070 43.785 ;
    RECT 0 43.855 0.070 44.205 ;
    RECT 0 44.275 0.070 44.625 ;
    RECT 0 44.695 0.070 45.045 ;
    RECT 0 45.115 0.070 45.465 ;
    RECT 0 45.535 0.070 45.885 ;
    RECT 0 45.955 0.070 46.305 ;
    RECT 0 46.375 0.070 46.725 ;
    RECT 0 46.795 0.070 47.145 ;
    RECT 0 47.215 0.070 47.565 ;
    RECT 0 47.635 0.070 47.985 ;
    RECT 0 48.055 0.070 48.405 ;
    RECT 0 48.475 0.070 48.825 ;
    RECT 0 48.895 0.070 49.245 ;
    RECT 0 49.315 0.070 49.665 ;
    RECT 0 49.735 0.070 50.085 ;
    RECT 0 50.155 0.070 50.505 ;
    RECT 0 50.575 0.070 50.925 ;
    RECT 0 50.995 0.070 51.345 ;
    RECT 0 51.415 0.070 51.765 ;
    RECT 0 51.835 0.070 52.185 ;
    RECT 0 52.255 0.070 52.605 ;
    RECT 0 52.675 0.070 53.025 ;
    RECT 0 53.095 0.070 53.445 ;
    RECT 0 53.515 0.070 53.865 ;
    RECT 0 53.935 0.070 54.285 ;
    RECT 0 54.355 0.070 54.705 ;
    RECT 0 54.775 0.070 55.125 ;
    RECT 0 55.195 0.070 55.545 ;
    RECT 0 55.615 0.070 55.965 ;
    RECT 0 56.035 0.070 56.385 ;
    RECT 0 56.455 0.070 56.805 ;
    RECT 0 56.875 0.070 57.225 ;
    RECT 0 57.295 0.070 57.645 ;
    RECT 0 57.715 0.070 58.065 ;
    RECT 0 58.135 0.070 58.485 ;
    RECT 0 58.555 0.070 58.905 ;
    RECT 0 58.975 0.070 59.325 ;
    RECT 0 59.395 0.070 59.745 ;
    RECT 0 59.815 0.070 60.165 ;
    RECT 0 60.235 0.070 60.585 ;
    RECT 0 60.655 0.070 61.005 ;
    RECT 0 61.075 0.070 61.425 ;
    RECT 0 61.495 0.070 61.845 ;
    RECT 0 61.915 0.070 62.265 ;
    RECT 0 62.335 0.070 62.685 ;
    RECT 0 62.755 0.070 63.105 ;
    RECT 0 63.175 0.070 63.525 ;
    RECT 0 63.595 0.070 63.945 ;
    RECT 0 64.015 0.070 64.365 ;
    RECT 0 64.435 0.070 64.785 ;
    RECT 0 64.855 0.070 65.205 ;
    RECT 0 65.275 0.070 65.625 ;
    RECT 0 65.695 0.070 66.045 ;
    RECT 0 66.115 0.070 66.465 ;
    RECT 0 66.535 0.070 66.885 ;
    RECT 0 66.955 0.070 67.305 ;
    RECT 0 67.375 0.070 67.725 ;
    RECT 0 67.795 0.070 68.145 ;
    RECT 0 68.215 0.070 68.565 ;
    RECT 0 68.635 0.070 68.985 ;
    RECT 0 69.055 0.070 69.405 ;
    RECT 0 69.475 0.070 69.825 ;
    RECT 0 69.895 0.070 70.245 ;
    RECT 0 70.315 0.070 70.665 ;
    RECT 0 70.735 0.070 71.085 ;
    RECT 0 71.155 0.070 71.505 ;
    RECT 0 71.575 0.070 71.925 ;
    RECT 0 71.995 0.070 72.345 ;
    RECT 0 72.415 0.070 72.765 ;
    RECT 0 72.835 0.070 73.185 ;
    RECT 0 73.255 0.070 73.605 ;
    RECT 0 73.675 0.070 74.025 ;
    RECT 0 74.095 0.070 74.445 ;
    RECT 0 74.515 0.070 74.865 ;
    RECT 0 74.935 0.070 75.285 ;
    RECT 0 75.355 0.070 75.705 ;
    RECT 0 75.775 0.070 76.125 ;
    RECT 0 76.195 0.070 76.545 ;
    RECT 0 76.615 0.070 76.965 ;
    RECT 0 77.035 0.070 77.385 ;
    RECT 0 77.455 0.070 77.805 ;
    RECT 0 77.875 0.070 78.225 ;
    RECT 0 78.295 0.070 78.645 ;
    RECT 0 78.715 0.070 79.065 ;
    RECT 0 79.135 0.070 79.485 ;
    RECT 0 79.555 0.070 79.905 ;
    RECT 0 79.975 0.070 80.325 ;
    RECT 0 80.395 0.070 80.745 ;
    RECT 0 80.815 0.070 81.165 ;
    RECT 0 81.235 0.070 81.585 ;
    RECT 0 81.655 0.070 82.005 ;
    RECT 0 82.075 0.070 82.425 ;
    RECT 0 82.495 0.070 82.845 ;
    RECT 0 82.915 0.070 83.265 ;
    RECT 0 83.335 0.070 83.685 ;
    RECT 0 83.755 0.070 84.105 ;
    RECT 0 84.175 0.070 84.525 ;
    RECT 0 84.595 0.070 84.945 ;
    RECT 0 85.015 0.070 85.365 ;
    RECT 0 85.435 0.070 85.785 ;
    RECT 0 85.855 0.070 86.205 ;
    RECT 0 86.275 0.070 86.625 ;
    RECT 0 86.695 0.070 87.045 ;
    RECT 0 87.115 0.070 87.465 ;
    RECT 0 87.535 0.070 87.885 ;
    RECT 0 87.955 0.070 88.305 ;
    RECT 0 88.375 0.070 88.725 ;
    RECT 0 88.795 0.070 89.145 ;
    RECT 0 89.215 0.070 89.565 ;
    RECT 0 89.635 0.070 89.985 ;
    RECT 0 90.055 0.070 90.405 ;
    RECT 0 90.475 0.070 90.825 ;
    RECT 0 90.895 0.070 91.245 ;
    RECT 0 91.315 0.070 91.665 ;
    RECT 0 91.735 0.070 92.085 ;
    RECT 0 92.155 0.070 92.505 ;
    RECT 0 92.575 0.070 92.925 ;
    RECT 0 92.995 0.070 93.345 ;
    RECT 0 93.415 0.070 93.765 ;
    RECT 0 93.835 0.070 94.185 ;
    RECT 0 94.255 0.070 94.605 ;
    RECT 0 94.675 0.070 95.025 ;
    RECT 0 95.095 0.070 95.445 ;
    RECT 0 95.515 0.070 95.865 ;
    RECT 0 95.935 0.070 96.285 ;
    RECT 0 96.355 0.070 96.705 ;
    RECT 0 96.775 0.070 97.125 ;
    RECT 0 97.195 0.070 97.545 ;
    RECT 0 97.615 0.070 97.965 ;
    RECT 0 98.035 0.070 98.385 ;
    RECT 0 98.455 0.070 98.805 ;
    RECT 0 98.875 0.070 99.225 ;
    RECT 0 99.295 0.070 99.645 ;
    RECT 0 99.715 0.070 100.065 ;
    RECT 0 100.135 0.070 100.485 ;
    RECT 0 100.555 0.070 100.905 ;
    RECT 0 100.975 0.070 101.325 ;
    RECT 0 101.395 0.070 101.745 ;
    RECT 0 101.815 0.070 102.165 ;
    RECT 0 102.235 0.070 102.585 ;
    RECT 0 102.655 0.070 103.005 ;
    RECT 0 103.075 0.070 103.425 ;
    RECT 0 103.495 0.070 103.845 ;
    RECT 0 103.915 0.070 104.265 ;
    RECT 0 104.335 0.070 104.685 ;
    RECT 0 104.755 0.070 105.105 ;
    RECT 0 105.175 0.070 105.525 ;
    RECT 0 105.595 0.070 105.945 ;
    RECT 0 106.015 0.070 106.365 ;
    RECT 0 106.435 0.070 106.785 ;
    RECT 0 106.855 0.070 107.205 ;
    RECT 0 107.275 0.070 107.625 ;
    RECT 0 107.695 0.070 108.045 ;
    RECT 0 108.115 0.070 108.465 ;
    RECT 0 108.535 0.070 108.885 ;
    RECT 0 108.955 0.070 109.305 ;
    RECT 0 109.375 0.070 109.725 ;
    RECT 0 109.795 0.070 110.145 ;
    RECT 0 110.215 0.070 110.565 ;
    RECT 0 110.635 0.070 110.985 ;
    RECT 0 111.055 0.070 111.405 ;
    RECT 0 111.475 0.070 111.825 ;
    RECT 0 111.895 0.070 112.245 ;
    RECT 0 112.315 0.070 112.665 ;
    RECT 0 112.735 0.070 113.085 ;
    RECT 0 113.155 0.070 113.505 ;
    RECT 0 113.575 0.070 113.925 ;
    RECT 0 113.995 0.070 114.345 ;
    RECT 0 114.415 0.070 114.765 ;
    RECT 0 114.835 0.070 115.185 ;
    RECT 0 115.255 0.070 115.605 ;
    RECT 0 115.675 0.070 116.025 ;
    RECT 0 116.095 0.070 116.445 ;
    RECT 0 116.515 0.070 116.865 ;
    RECT 0 116.935 0.070 117.285 ;
    RECT 0 117.355 0.070 117.705 ;
    RECT 0 117.775 0.070 118.125 ;
    RECT 0 118.195 0.070 118.545 ;
    RECT 0 118.615 0.070 118.965 ;
    RECT 0 119.035 0.070 119.385 ;
    RECT 0 119.455 0.070 119.805 ;
    RECT 0 119.875 0.070 120.225 ;
    RECT 0 120.295 0.070 120.645 ;
    RECT 0 120.715 0.070 121.065 ;
    RECT 0 121.135 0.070 121.485 ;
    RECT 0 121.555 0.070 121.905 ;
    RECT 0 121.975 0.070 122.325 ;
    RECT 0 122.395 0.070 122.745 ;
    RECT 0 122.815 0.070 123.165 ;
    RECT 0 123.235 0.070 123.585 ;
    RECT 0 123.655 0.070 124.005 ;
    RECT 0 124.075 0.070 124.425 ;
    RECT 0 124.495 0.070 124.845 ;
    RECT 0 124.915 0.070 125.265 ;
    RECT 0 125.335 0.070 125.685 ;
    RECT 0 125.755 0.070 126.105 ;
    RECT 0 126.175 0.070 126.525 ;
    RECT 0 126.595 0.070 126.945 ;
    RECT 0 127.015 0.070 127.365 ;
    RECT 0 127.435 0.070 127.785 ;
    RECT 0 127.855 0.070 128.205 ;
    RECT 0 128.275 0.070 128.625 ;
    RECT 0 128.695 0.070 129.045 ;
    RECT 0 129.115 0.070 129.465 ;
    RECT 0 129.535 0.070 129.885 ;
    RECT 0 129.955 0.070 130.305 ;
    RECT 0 130.375 0.070 130.725 ;
    RECT 0 130.795 0.070 131.145 ;
    RECT 0 131.215 0.070 131.565 ;
    RECT 0 131.635 0.070 131.985 ;
    RECT 0 132.055 0.070 132.405 ;
    RECT 0 132.475 0.070 132.825 ;
    RECT 0 132.895 0.070 133.245 ;
    RECT 0 133.315 0.070 133.665 ;
    RECT 0 133.735 0.070 134.085 ;
    RECT 0 134.155 0.070 134.505 ;
    RECT 0 134.575 0.070 134.925 ;
    RECT 0 134.995 0.070 135.345 ;
    RECT 0 135.415 0.070 135.765 ;
    RECT 0 135.835 0.070 136.185 ;
    RECT 0 136.255 0.070 136.605 ;
    RECT 0 136.675 0.070 137.025 ;
    RECT 0 137.095 0.070 137.445 ;
    RECT 0 137.515 0.070 137.865 ;
    RECT 0 137.935 0.070 138.285 ;
    RECT 0 138.355 0.070 138.705 ;
    RECT 0 138.775 0.070 139.125 ;
    RECT 0 139.195 0.070 139.545 ;
    RECT 0 139.615 0.070 139.965 ;
    RECT 0 140.035 0.070 140.385 ;
    RECT 0 140.455 0.070 140.805 ;
    RECT 0 140.875 0.070 141.225 ;
    RECT 0 141.295 0.070 141.645 ;
    RECT 0 141.715 0.070 142.065 ;
    RECT 0 142.135 0.070 142.485 ;
    RECT 0 142.555 0.070 142.905 ;
    RECT 0 142.975 0.070 143.325 ;
    RECT 0 143.395 0.070 143.745 ;
    RECT 0 143.815 0.070 144.165 ;
    RECT 0 144.235 0.070 144.585 ;
    RECT 0 144.655 0.070 145.005 ;
    RECT 0 145.075 0.070 145.425 ;
    RECT 0 145.495 0.070 145.845 ;
    RECT 0 145.915 0.070 146.265 ;
    RECT 0 146.335 0.070 146.685 ;
    RECT 0 146.755 0.070 147.105 ;
    RECT 0 147.175 0.070 147.525 ;
    RECT 0 147.595 0.070 147.945 ;
    RECT 0 148.015 0.070 148.365 ;
    RECT 0 148.435 0.070 148.785 ;
    RECT 0 148.855 0.070 149.205 ;
    RECT 0 149.275 0.070 149.625 ;
    RECT 0 149.695 0.070 150.045 ;
    RECT 0 150.115 0.070 150.465 ;
    RECT 0 150.535 0.070 150.885 ;
    RECT 0 150.955 0.070 151.305 ;
    RECT 0 151.375 0.070 151.725 ;
    RECT 0 151.795 0.070 152.145 ;
    RECT 0 152.215 0.070 152.565 ;
    RECT 0 152.635 0.070 152.985 ;
    RECT 0 153.055 0.070 153.405 ;
    RECT 0 153.475 0.070 153.825 ;
    RECT 0 153.895 0.070 154.245 ;
    RECT 0 154.315 0.070 154.665 ;
    RECT 0 154.735 0.070 155.085 ;
    RECT 0 155.155 0.070 155.505 ;
    RECT 0 155.575 0.070 155.925 ;
    RECT 0 155.995 0.070 156.345 ;
    RECT 0 156.415 0.070 156.765 ;
    RECT 0 156.835 0.070 157.185 ;
    RECT 0 157.255 0.070 157.605 ;
    RECT 0 157.675 0.070 158.025 ;
    RECT 0 158.095 0.070 158.445 ;
    RECT 0 158.515 0.070 158.865 ;
    RECT 0 158.935 0.070 159.285 ;
    RECT 0 159.355 0.070 159.705 ;
    RECT 0 159.775 0.070 160.125 ;
    RECT 0 160.195 0.070 160.545 ;
    RECT 0 160.615 0.070 160.965 ;
    RECT 0 161.035 0.070 161.385 ;
    RECT 0 161.455 0.070 161.805 ;
    RECT 0 161.875 0.070 162.225 ;
    RECT 0 162.295 0.070 162.645 ;
    RECT 0 162.715 0.070 163.065 ;
    RECT 0 163.135 0.070 163.485 ;
    RECT 0 163.555 0.070 163.905 ;
    RECT 0 163.975 0.070 164.325 ;
    RECT 0 164.395 0.070 164.745 ;
    RECT 0 164.815 0.070 165.165 ;
    RECT 0 165.235 0.070 165.585 ;
    RECT 0 165.655 0.070 166.005 ;
    RECT 0 166.075 0.070 166.425 ;
    RECT 0 166.495 0.070 166.845 ;
    RECT 0 166.915 0.070 167.265 ;
    RECT 0 167.335 0.070 167.685 ;
    RECT 0 167.755 0.070 168.105 ;
    RECT 0 168.175 0.070 168.525 ;
    RECT 0 168.595 0.070 168.945 ;
    RECT 0 169.015 0.070 169.365 ;
    RECT 0 169.435 0.070 169.785 ;
    RECT 0 169.855 0.070 170.205 ;
    RECT 0 170.275 0.070 170.625 ;
    RECT 0 170.695 0.070 171.045 ;
    RECT 0 171.115 0.070 171.465 ;
    RECT 0 171.535 0.070 171.885 ;
    RECT 0 171.955 0.070 172.305 ;
    RECT 0 172.375 0.070 172.725 ;
    RECT 0 172.795 0.070 173.145 ;
    RECT 0 173.215 0.070 173.565 ;
    RECT 0 173.635 0.070 173.985 ;
    RECT 0 174.055 0.070 174.405 ;
    RECT 0 174.475 0.070 174.825 ;
    RECT 0 174.895 0.070 175.245 ;
    RECT 0 175.315 0.070 175.665 ;
    RECT 0 175.735 0.070 176.085 ;
    RECT 0 176.155 0.070 176.505 ;
    RECT 0 176.575 0.070 176.925 ;
    RECT 0 176.995 0.070 177.345 ;
    RECT 0 177.415 0.070 177.765 ;
    RECT 0 177.835 0.070 178.185 ;
    RECT 0 178.255 0.070 178.605 ;
    RECT 0 178.675 0.070 179.025 ;
    RECT 0 179.095 0.070 179.445 ;
    RECT 0 179.515 0.070 179.865 ;
    RECT 0 179.935 0.070 180.285 ;
    RECT 0 180.355 0.070 180.705 ;
    RECT 0 180.775 0.070 181.125 ;
    RECT 0 181.195 0.070 181.545 ;
    RECT 0 181.615 0.070 181.965 ;
    RECT 0 182.035 0.070 182.385 ;
    RECT 0 182.455 0.070 182.805 ;
    RECT 0 182.875 0.070 183.225 ;
    RECT 0 183.295 0.070 183.645 ;
    RECT 0 183.715 0.070 184.065 ;
    RECT 0 184.135 0.070 184.485 ;
    RECT 0 184.555 0.070 184.905 ;
    RECT 0 184.975 0.070 185.325 ;
    RECT 0 185.395 0.070 185.745 ;
    RECT 0 185.815 0.070 186.165 ;
    RECT 0 186.235 0.070 186.585 ;
    RECT 0 186.655 0.070 187.005 ;
    RECT 0 187.075 0.070 187.425 ;
    RECT 0 187.495 0.070 187.845 ;
    RECT 0 187.915 0.070 188.265 ;
    RECT 0 188.335 0.070 188.685 ;
    RECT 0 188.755 0.070 189.105 ;
    RECT 0 189.175 0.070 189.525 ;
    RECT 0 189.595 0.070 189.945 ;
    RECT 0 190.015 0.070 190.365 ;
    RECT 0 190.435 0.070 190.785 ;
    RECT 0 190.855 0.070 191.205 ;
    RECT 0 191.275 0.070 191.625 ;
    RECT 0 191.695 0.070 192.045 ;
    RECT 0 192.115 0.070 192.465 ;
    RECT 0 192.535 0.070 192.885 ;
    RECT 0 192.955 0.070 193.305 ;
    RECT 0 193.375 0.070 193.725 ;
    RECT 0 193.795 0.070 194.145 ;
    RECT 0 194.215 0.070 194.565 ;
    RECT 0 194.635 0.070 194.985 ;
    RECT 0 195.055 0.070 195.405 ;
    RECT 0 195.475 0.070 195.825 ;
    RECT 0 195.895 0.070 196.245 ;
    RECT 0 196.315 0.070 196.665 ;
    RECT 0 196.735 0.070 197.085 ;
    RECT 0 197.155 0.070 197.505 ;
    RECT 0 197.575 0.070 197.925 ;
    RECT 0 197.995 0.070 198.345 ;
    RECT 0 198.415 0.070 198.765 ;
    RECT 0 198.835 0.070 199.185 ;
    RECT 0 199.255 0.070 199.605 ;
    RECT 0 199.675 0.070 200.025 ;
    RECT 0 200.095 0.070 200.445 ;
    RECT 0 200.515 0.070 200.865 ;
    RECT 0 200.935 0.070 201.285 ;
    RECT 0 201.355 0.070 201.705 ;
    RECT 0 201.775 0.070 202.125 ;
    RECT 0 202.195 0.070 202.545 ;
    RECT 0 202.615 0.070 202.965 ;
    RECT 0 203.035 0.070 203.385 ;
    RECT 0 203.455 0.070 203.805 ;
    RECT 0 203.875 0.070 204.225 ;
    RECT 0 204.295 0.070 204.645 ;
    RECT 0 204.715 0.070 205.065 ;
    RECT 0 205.135 0.070 205.485 ;
    RECT 0 205.555 0.070 205.905 ;
    RECT 0 205.975 0.070 206.325 ;
    RECT 0 206.395 0.070 206.745 ;
    RECT 0 206.815 0.070 207.165 ;
    RECT 0 207.235 0.070 207.585 ;
    RECT 0 207.655 0.070 208.005 ;
    RECT 0 208.075 0.070 208.425 ;
    RECT 0 208.495 0.070 208.845 ;
    RECT 0 208.915 0.070 209.265 ;
    RECT 0 209.335 0.070 209.685 ;
    RECT 0 209.755 0.070 210.105 ;
    RECT 0 210.175 0.070 210.525 ;
    RECT 0 210.595 0.070 210.945 ;
    RECT 0 211.015 0.070 211.365 ;
    RECT 0 211.435 0.070 211.785 ;
    RECT 0 211.855 0.070 212.205 ;
    RECT 0 212.275 0.070 212.625 ;
    RECT 0 212.695 0.070 213.045 ;
    RECT 0 213.115 0.070 213.465 ;
    RECT 0 213.535 0.070 213.885 ;
    RECT 0 213.955 0.070 214.305 ;
    RECT 0 214.375 0.070 214.725 ;
    RECT 0 214.795 0.070 215.145 ;
    RECT 0 215.215 0.070 215.565 ;
    RECT 0 215.635 0.070 215.985 ;
    RECT 0 216.055 0.070 244.545 ;
    RECT 0 244.615 0.070 244.965 ;
    RECT 0 245.035 0.070 245.385 ;
    RECT 0 245.455 0.070 245.805 ;
    RECT 0 245.875 0.070 246.225 ;
    RECT 0 246.295 0.070 246.645 ;
    RECT 0 246.715 0.070 247.065 ;
    RECT 0 247.135 0.070 247.485 ;
    RECT 0 247.555 0.070 247.905 ;
    RECT 0 247.975 0.070 248.325 ;
    RECT 0 248.395 0.070 248.745 ;
    RECT 0 248.815 0.070 249.165 ;
    RECT 0 249.235 0.070 249.585 ;
    RECT 0 249.655 0.070 250.005 ;
    RECT 0 250.075 0.070 250.425 ;
    RECT 0 250.495 0.070 250.845 ;
    RECT 0 250.915 0.070 251.265 ;
    RECT 0 251.335 0.070 251.685 ;
    RECT 0 251.755 0.070 252.105 ;
    RECT 0 252.175 0.070 252.525 ;
    RECT 0 252.595 0.070 252.945 ;
    RECT 0 253.015 0.070 253.365 ;
    RECT 0 253.435 0.070 253.785 ;
    RECT 0 253.855 0.070 254.205 ;
    RECT 0 254.275 0.070 254.625 ;
    RECT 0 254.695 0.070 255.045 ;
    RECT 0 255.115 0.070 255.465 ;
    RECT 0 255.535 0.070 255.885 ;
    RECT 0 255.955 0.070 256.305 ;
    RECT 0 256.375 0.070 256.725 ;
    RECT 0 256.795 0.070 257.145 ;
    RECT 0 257.215 0.070 257.565 ;
    RECT 0 257.635 0.070 257.985 ;
    RECT 0 258.055 0.070 258.405 ;
    RECT 0 258.475 0.070 258.825 ;
    RECT 0 258.895 0.070 259.245 ;
    RECT 0 259.315 0.070 259.665 ;
    RECT 0 259.735 0.070 260.085 ;
    RECT 0 260.155 0.070 260.505 ;
    RECT 0 260.575 0.070 260.925 ;
    RECT 0 260.995 0.070 261.345 ;
    RECT 0 261.415 0.070 261.765 ;
    RECT 0 261.835 0.070 262.185 ;
    RECT 0 262.255 0.070 262.605 ;
    RECT 0 262.675 0.070 263.025 ;
    RECT 0 263.095 0.070 263.445 ;
    RECT 0 263.515 0.070 263.865 ;
    RECT 0 263.935 0.070 264.285 ;
    RECT 0 264.355 0.070 264.705 ;
    RECT 0 264.775 0.070 265.125 ;
    RECT 0 265.195 0.070 265.545 ;
    RECT 0 265.615 0.070 265.965 ;
    RECT 0 266.035 0.070 266.385 ;
    RECT 0 266.455 0.070 266.805 ;
    RECT 0 266.875 0.070 267.225 ;
    RECT 0 267.295 0.070 267.645 ;
    RECT 0 267.715 0.070 268.065 ;
    RECT 0 268.135 0.070 268.485 ;
    RECT 0 268.555 0.070 268.905 ;
    RECT 0 268.975 0.070 269.325 ;
    RECT 0 269.395 0.070 269.745 ;
    RECT 0 269.815 0.070 270.165 ;
    RECT 0 270.235 0.070 270.585 ;
    RECT 0 270.655 0.070 271.005 ;
    RECT 0 271.075 0.070 271.425 ;
    RECT 0 271.495 0.070 271.845 ;
    RECT 0 271.915 0.070 272.265 ;
    RECT 0 272.335 0.070 272.685 ;
    RECT 0 272.755 0.070 273.105 ;
    RECT 0 273.175 0.070 273.525 ;
    RECT 0 273.595 0.070 273.945 ;
    RECT 0 274.015 0.070 274.365 ;
    RECT 0 274.435 0.070 274.785 ;
    RECT 0 274.855 0.070 275.205 ;
    RECT 0 275.275 0.070 275.625 ;
    RECT 0 275.695 0.070 276.045 ;
    RECT 0 276.115 0.070 276.465 ;
    RECT 0 276.535 0.070 276.885 ;
    RECT 0 276.955 0.070 277.305 ;
    RECT 0 277.375 0.070 277.725 ;
    RECT 0 277.795 0.070 278.145 ;
    RECT 0 278.215 0.070 278.565 ;
    RECT 0 278.635 0.070 278.985 ;
    RECT 0 279.055 0.070 279.405 ;
    RECT 0 279.475 0.070 279.825 ;
    RECT 0 279.895 0.070 280.245 ;
    RECT 0 280.315 0.070 280.665 ;
    RECT 0 280.735 0.070 281.085 ;
    RECT 0 281.155 0.070 281.505 ;
    RECT 0 281.575 0.070 281.925 ;
    RECT 0 281.995 0.070 282.345 ;
    RECT 0 282.415 0.070 282.765 ;
    RECT 0 282.835 0.070 283.185 ;
    RECT 0 283.255 0.070 283.605 ;
    RECT 0 283.675 0.070 284.025 ;
    RECT 0 284.095 0.070 284.445 ;
    RECT 0 284.515 0.070 284.865 ;
    RECT 0 284.935 0.070 285.285 ;
    RECT 0 285.355 0.070 285.705 ;
    RECT 0 285.775 0.070 286.125 ;
    RECT 0 286.195 0.070 286.545 ;
    RECT 0 286.615 0.070 286.965 ;
    RECT 0 287.035 0.070 287.385 ;
    RECT 0 287.455 0.070 287.805 ;
    RECT 0 287.875 0.070 288.225 ;
    RECT 0 288.295 0.070 288.645 ;
    RECT 0 288.715 0.070 289.065 ;
    RECT 0 289.135 0.070 289.485 ;
    RECT 0 289.555 0.070 289.905 ;
    RECT 0 289.975 0.070 290.325 ;
    RECT 0 290.395 0.070 290.745 ;
    RECT 0 290.815 0.070 291.165 ;
    RECT 0 291.235 0.070 291.585 ;
    RECT 0 291.655 0.070 292.005 ;
    RECT 0 292.075 0.070 292.425 ;
    RECT 0 292.495 0.070 292.845 ;
    RECT 0 292.915 0.070 293.265 ;
    RECT 0 293.335 0.070 293.685 ;
    RECT 0 293.755 0.070 294.105 ;
    RECT 0 294.175 0.070 294.525 ;
    RECT 0 294.595 0.070 294.945 ;
    RECT 0 295.015 0.070 295.365 ;
    RECT 0 295.435 0.070 295.785 ;
    RECT 0 295.855 0.070 296.205 ;
    RECT 0 296.275 0.070 296.625 ;
    RECT 0 296.695 0.070 297.045 ;
    RECT 0 297.115 0.070 297.465 ;
    RECT 0 297.535 0.070 297.885 ;
    RECT 0 297.955 0.070 298.305 ;
    RECT 0 298.375 0.070 298.725 ;
    RECT 0 298.795 0.070 299.145 ;
    RECT 0 299.215 0.070 299.565 ;
    RECT 0 299.635 0.070 299.985 ;
    RECT 0 300.055 0.070 300.405 ;
    RECT 0 300.475 0.070 300.825 ;
    RECT 0 300.895 0.070 301.245 ;
    RECT 0 301.315 0.070 301.665 ;
    RECT 0 301.735 0.070 302.085 ;
    RECT 0 302.155 0.070 302.505 ;
    RECT 0 302.575 0.070 302.925 ;
    RECT 0 302.995 0.070 303.345 ;
    RECT 0 303.415 0.070 303.765 ;
    RECT 0 303.835 0.070 304.185 ;
    RECT 0 304.255 0.070 304.605 ;
    RECT 0 304.675 0.070 305.025 ;
    RECT 0 305.095 0.070 305.445 ;
    RECT 0 305.515 0.070 305.865 ;
    RECT 0 305.935 0.070 306.285 ;
    RECT 0 306.355 0.070 306.705 ;
    RECT 0 306.775 0.070 307.125 ;
    RECT 0 307.195 0.070 307.545 ;
    RECT 0 307.615 0.070 307.965 ;
    RECT 0 308.035 0.070 308.385 ;
    RECT 0 308.455 0.070 308.805 ;
    RECT 0 308.875 0.070 309.225 ;
    RECT 0 309.295 0.070 309.645 ;
    RECT 0 309.715 0.070 310.065 ;
    RECT 0 310.135 0.070 310.485 ;
    RECT 0 310.555 0.070 310.905 ;
    RECT 0 310.975 0.070 311.325 ;
    RECT 0 311.395 0.070 311.745 ;
    RECT 0 311.815 0.070 312.165 ;
    RECT 0 312.235 0.070 312.585 ;
    RECT 0 312.655 0.070 313.005 ;
    RECT 0 313.075 0.070 313.425 ;
    RECT 0 313.495 0.070 313.845 ;
    RECT 0 313.915 0.070 314.265 ;
    RECT 0 314.335 0.070 314.685 ;
    RECT 0 314.755 0.070 315.105 ;
    RECT 0 315.175 0.070 315.525 ;
    RECT 0 315.595 0.070 315.945 ;
    RECT 0 316.015 0.070 316.365 ;
    RECT 0 316.435 0.070 316.785 ;
    RECT 0 316.855 0.070 317.205 ;
    RECT 0 317.275 0.070 317.625 ;
    RECT 0 317.695 0.070 318.045 ;
    RECT 0 318.115 0.070 318.465 ;
    RECT 0 318.535 0.070 318.885 ;
    RECT 0 318.955 0.070 319.305 ;
    RECT 0 319.375 0.070 319.725 ;
    RECT 0 319.795 0.070 320.145 ;
    RECT 0 320.215 0.070 320.565 ;
    RECT 0 320.635 0.070 320.985 ;
    RECT 0 321.055 0.070 321.405 ;
    RECT 0 321.475 0.070 321.825 ;
    RECT 0 321.895 0.070 322.245 ;
    RECT 0 322.315 0.070 322.665 ;
    RECT 0 322.735 0.070 323.085 ;
    RECT 0 323.155 0.070 323.505 ;
    RECT 0 323.575 0.070 323.925 ;
    RECT 0 323.995 0.070 324.345 ;
    RECT 0 324.415 0.070 324.765 ;
    RECT 0 324.835 0.070 325.185 ;
    RECT 0 325.255 0.070 325.605 ;
    RECT 0 325.675 0.070 326.025 ;
    RECT 0 326.095 0.070 326.445 ;
    RECT 0 326.515 0.070 326.865 ;
    RECT 0 326.935 0.070 327.285 ;
    RECT 0 327.355 0.070 327.705 ;
    RECT 0 327.775 0.070 328.125 ;
    RECT 0 328.195 0.070 328.545 ;
    RECT 0 328.615 0.070 328.965 ;
    RECT 0 329.035 0.070 329.385 ;
    RECT 0 329.455 0.070 329.805 ;
    RECT 0 329.875 0.070 330.225 ;
    RECT 0 330.295 0.070 330.645 ;
    RECT 0 330.715 0.070 331.065 ;
    RECT 0 331.135 0.070 331.485 ;
    RECT 0 331.555 0.070 331.905 ;
    RECT 0 331.975 0.070 332.325 ;
    RECT 0 332.395 0.070 332.745 ;
    RECT 0 332.815 0.070 333.165 ;
    RECT 0 333.235 0.070 333.585 ;
    RECT 0 333.655 0.070 334.005 ;
    RECT 0 334.075 0.070 334.425 ;
    RECT 0 334.495 0.070 334.845 ;
    RECT 0 334.915 0.070 335.265 ;
    RECT 0 335.335 0.070 335.685 ;
    RECT 0 335.755 0.070 336.105 ;
    RECT 0 336.175 0.070 336.525 ;
    RECT 0 336.595 0.070 336.945 ;
    RECT 0 337.015 0.070 337.365 ;
    RECT 0 337.435 0.070 337.785 ;
    RECT 0 337.855 0.070 338.205 ;
    RECT 0 338.275 0.070 338.625 ;
    RECT 0 338.695 0.070 339.045 ;
    RECT 0 339.115 0.070 339.465 ;
    RECT 0 339.535 0.070 339.885 ;
    RECT 0 339.955 0.070 340.305 ;
    RECT 0 340.375 0.070 340.725 ;
    RECT 0 340.795 0.070 341.145 ;
    RECT 0 341.215 0.070 341.565 ;
    RECT 0 341.635 0.070 341.985 ;
    RECT 0 342.055 0.070 342.405 ;
    RECT 0 342.475 0.070 342.825 ;
    RECT 0 342.895 0.070 343.245 ;
    RECT 0 343.315 0.070 343.665 ;
    RECT 0 343.735 0.070 344.085 ;
    RECT 0 344.155 0.070 344.505 ;
    RECT 0 344.575 0.070 344.925 ;
    RECT 0 344.995 0.070 345.345 ;
    RECT 0 345.415 0.070 345.765 ;
    RECT 0 345.835 0.070 346.185 ;
    RECT 0 346.255 0.070 346.605 ;
    RECT 0 346.675 0.070 347.025 ;
    RECT 0 347.095 0.070 347.445 ;
    RECT 0 347.515 0.070 347.865 ;
    RECT 0 347.935 0.070 348.285 ;
    RECT 0 348.355 0.070 348.705 ;
    RECT 0 348.775 0.070 349.125 ;
    RECT 0 349.195 0.070 349.545 ;
    RECT 0 349.615 0.070 349.965 ;
    RECT 0 350.035 0.070 350.385 ;
    RECT 0 350.455 0.070 350.805 ;
    RECT 0 350.875 0.070 351.225 ;
    RECT 0 351.295 0.070 351.645 ;
    RECT 0 351.715 0.070 352.065 ;
    RECT 0 352.135 0.070 352.485 ;
    RECT 0 352.555 0.070 352.905 ;
    RECT 0 352.975 0.070 353.325 ;
    RECT 0 353.395 0.070 353.745 ;
    RECT 0 353.815 0.070 354.165 ;
    RECT 0 354.235 0.070 354.585 ;
    RECT 0 354.655 0.070 355.005 ;
    RECT 0 355.075 0.070 355.425 ;
    RECT 0 355.495 0.070 355.845 ;
    RECT 0 355.915 0.070 356.265 ;
    RECT 0 356.335 0.070 356.685 ;
    RECT 0 356.755 0.070 357.105 ;
    RECT 0 357.175 0.070 357.525 ;
    RECT 0 357.595 0.070 357.945 ;
    RECT 0 358.015 0.070 358.365 ;
    RECT 0 358.435 0.070 358.785 ;
    RECT 0 358.855 0.070 359.205 ;
    RECT 0 359.275 0.070 359.625 ;
    RECT 0 359.695 0.070 360.045 ;
    RECT 0 360.115 0.070 360.465 ;
    RECT 0 360.535 0.070 360.885 ;
    RECT 0 360.955 0.070 361.305 ;
    RECT 0 361.375 0.070 361.725 ;
    RECT 0 361.795 0.070 362.145 ;
    RECT 0 362.215 0.070 362.565 ;
    RECT 0 362.635 0.070 362.985 ;
    RECT 0 363.055 0.070 363.405 ;
    RECT 0 363.475 0.070 363.825 ;
    RECT 0 363.895 0.070 364.245 ;
    RECT 0 364.315 0.070 364.665 ;
    RECT 0 364.735 0.070 365.085 ;
    RECT 0 365.155 0.070 365.505 ;
    RECT 0 365.575 0.070 365.925 ;
    RECT 0 365.995 0.070 366.345 ;
    RECT 0 366.415 0.070 366.765 ;
    RECT 0 366.835 0.070 367.185 ;
    RECT 0 367.255 0.070 367.605 ;
    RECT 0 367.675 0.070 368.025 ;
    RECT 0 368.095 0.070 368.445 ;
    RECT 0 368.515 0.070 368.865 ;
    RECT 0 368.935 0.070 369.285 ;
    RECT 0 369.355 0.070 369.705 ;
    RECT 0 369.775 0.070 370.125 ;
    RECT 0 370.195 0.070 370.545 ;
    RECT 0 370.615 0.070 370.965 ;
    RECT 0 371.035 0.070 371.385 ;
    RECT 0 371.455 0.070 371.805 ;
    RECT 0 371.875 0.070 372.225 ;
    RECT 0 372.295 0.070 372.645 ;
    RECT 0 372.715 0.070 373.065 ;
    RECT 0 373.135 0.070 373.485 ;
    RECT 0 373.555 0.070 373.905 ;
    RECT 0 373.975 0.070 374.325 ;
    RECT 0 374.395 0.070 374.745 ;
    RECT 0 374.815 0.070 375.165 ;
    RECT 0 375.235 0.070 375.585 ;
    RECT 0 375.655 0.070 376.005 ;
    RECT 0 376.075 0.070 376.425 ;
    RECT 0 376.495 0.070 376.845 ;
    RECT 0 376.915 0.070 377.265 ;
    RECT 0 377.335 0.070 377.685 ;
    RECT 0 377.755 0.070 378.105 ;
    RECT 0 378.175 0.070 378.525 ;
    RECT 0 378.595 0.070 378.945 ;
    RECT 0 379.015 0.070 379.365 ;
    RECT 0 379.435 0.070 379.785 ;
    RECT 0 379.855 0.070 380.205 ;
    RECT 0 380.275 0.070 380.625 ;
    RECT 0 380.695 0.070 381.045 ;
    RECT 0 381.115 0.070 381.465 ;
    RECT 0 381.535 0.070 381.885 ;
    RECT 0 381.955 0.070 382.305 ;
    RECT 0 382.375 0.070 382.725 ;
    RECT 0 382.795 0.070 383.145 ;
    RECT 0 383.215 0.070 383.565 ;
    RECT 0 383.635 0.070 383.985 ;
    RECT 0 384.055 0.070 384.405 ;
    RECT 0 384.475 0.070 384.825 ;
    RECT 0 384.895 0.070 385.245 ;
    RECT 0 385.315 0.070 385.665 ;
    RECT 0 385.735 0.070 386.085 ;
    RECT 0 386.155 0.070 386.505 ;
    RECT 0 386.575 0.070 386.925 ;
    RECT 0 386.995 0.070 387.345 ;
    RECT 0 387.415 0.070 387.765 ;
    RECT 0 387.835 0.070 388.185 ;
    RECT 0 388.255 0.070 388.605 ;
    RECT 0 388.675 0.070 389.025 ;
    RECT 0 389.095 0.070 389.445 ;
    RECT 0 389.515 0.070 389.865 ;
    RECT 0 389.935 0.070 390.285 ;
    RECT 0 390.355 0.070 390.705 ;
    RECT 0 390.775 0.070 391.125 ;
    RECT 0 391.195 0.070 391.545 ;
    RECT 0 391.615 0.070 391.965 ;
    RECT 0 392.035 0.070 392.385 ;
    RECT 0 392.455 0.070 392.805 ;
    RECT 0 392.875 0.070 393.225 ;
    RECT 0 393.295 0.070 393.645 ;
    RECT 0 393.715 0.070 394.065 ;
    RECT 0 394.135 0.070 394.485 ;
    RECT 0 394.555 0.070 394.905 ;
    RECT 0 394.975 0.070 395.325 ;
    RECT 0 395.395 0.070 395.745 ;
    RECT 0 395.815 0.070 396.165 ;
    RECT 0 396.235 0.070 396.585 ;
    RECT 0 396.655 0.070 397.005 ;
    RECT 0 397.075 0.070 397.425 ;
    RECT 0 397.495 0.070 397.845 ;
    RECT 0 397.915 0.070 398.265 ;
    RECT 0 398.335 0.070 398.685 ;
    RECT 0 398.755 0.070 399.105 ;
    RECT 0 399.175 0.070 399.525 ;
    RECT 0 399.595 0.070 399.945 ;
    RECT 0 400.015 0.070 400.365 ;
    RECT 0 400.435 0.070 400.785 ;
    RECT 0 400.855 0.070 401.205 ;
    RECT 0 401.275 0.070 401.625 ;
    RECT 0 401.695 0.070 402.045 ;
    RECT 0 402.115 0.070 402.465 ;
    RECT 0 402.535 0.070 402.885 ;
    RECT 0 402.955 0.070 403.305 ;
    RECT 0 403.375 0.070 403.725 ;
    RECT 0 403.795 0.070 404.145 ;
    RECT 0 404.215 0.070 404.565 ;
    RECT 0 404.635 0.070 404.985 ;
    RECT 0 405.055 0.070 405.405 ;
    RECT 0 405.475 0.070 405.825 ;
    RECT 0 405.895 0.070 406.245 ;
    RECT 0 406.315 0.070 406.665 ;
    RECT 0 406.735 0.070 407.085 ;
    RECT 0 407.155 0.070 407.505 ;
    RECT 0 407.575 0.070 407.925 ;
    RECT 0 407.995 0.070 408.345 ;
    RECT 0 408.415 0.070 408.765 ;
    RECT 0 408.835 0.070 409.185 ;
    RECT 0 409.255 0.070 409.605 ;
    RECT 0 409.675 0.070 410.025 ;
    RECT 0 410.095 0.070 410.445 ;
    RECT 0 410.515 0.070 410.865 ;
    RECT 0 410.935 0.070 411.285 ;
    RECT 0 411.355 0.070 411.705 ;
    RECT 0 411.775 0.070 412.125 ;
    RECT 0 412.195 0.070 412.545 ;
    RECT 0 412.615 0.070 412.965 ;
    RECT 0 413.035 0.070 413.385 ;
    RECT 0 413.455 0.070 413.805 ;
    RECT 0 413.875 0.070 414.225 ;
    RECT 0 414.295 0.070 414.645 ;
    RECT 0 414.715 0.070 415.065 ;
    RECT 0 415.135 0.070 415.485 ;
    RECT 0 415.555 0.070 415.905 ;
    RECT 0 415.975 0.070 416.325 ;
    RECT 0 416.395 0.070 416.745 ;
    RECT 0 416.815 0.070 417.165 ;
    RECT 0 417.235 0.070 417.585 ;
    RECT 0 417.655 0.070 418.005 ;
    RECT 0 418.075 0.070 418.425 ;
    RECT 0 418.495 0.070 418.845 ;
    RECT 0 418.915 0.070 419.265 ;
    RECT 0 419.335 0.070 419.685 ;
    RECT 0 419.755 0.070 420.105 ;
    RECT 0 420.175 0.070 420.525 ;
    RECT 0 420.595 0.070 420.945 ;
    RECT 0 421.015 0.070 421.365 ;
    RECT 0 421.435 0.070 421.785 ;
    RECT 0 421.855 0.070 422.205 ;
    RECT 0 422.275 0.070 422.625 ;
    RECT 0 422.695 0.070 423.045 ;
    RECT 0 423.115 0.070 423.465 ;
    RECT 0 423.535 0.070 423.885 ;
    RECT 0 423.955 0.070 424.305 ;
    RECT 0 424.375 0.070 424.725 ;
    RECT 0 424.795 0.070 425.145 ;
    RECT 0 425.215 0.070 425.565 ;
    RECT 0 425.635 0.070 425.985 ;
    RECT 0 426.055 0.070 426.405 ;
    RECT 0 426.475 0.070 426.825 ;
    RECT 0 426.895 0.070 427.245 ;
    RECT 0 427.315 0.070 427.665 ;
    RECT 0 427.735 0.070 428.085 ;
    RECT 0 428.155 0.070 428.505 ;
    RECT 0 428.575 0.070 428.925 ;
    RECT 0 428.995 0.070 429.345 ;
    RECT 0 429.415 0.070 429.765 ;
    RECT 0 429.835 0.070 430.185 ;
    RECT 0 430.255 0.070 430.605 ;
    RECT 0 430.675 0.070 431.025 ;
    RECT 0 431.095 0.070 431.445 ;
    RECT 0 431.515 0.070 431.865 ;
    RECT 0 431.935 0.070 432.285 ;
    RECT 0 432.355 0.070 432.705 ;
    RECT 0 432.775 0.070 433.125 ;
    RECT 0 433.195 0.070 433.545 ;
    RECT 0 433.615 0.070 433.965 ;
    RECT 0 434.035 0.070 434.385 ;
    RECT 0 434.455 0.070 434.805 ;
    RECT 0 434.875 0.070 435.225 ;
    RECT 0 435.295 0.070 435.645 ;
    RECT 0 435.715 0.070 436.065 ;
    RECT 0 436.135 0.070 436.485 ;
    RECT 0 436.555 0.070 436.905 ;
    RECT 0 436.975 0.070 437.325 ;
    RECT 0 437.395 0.070 437.745 ;
    RECT 0 437.815 0.070 438.165 ;
    RECT 0 438.235 0.070 438.585 ;
    RECT 0 438.655 0.070 439.005 ;
    RECT 0 439.075 0.070 439.425 ;
    RECT 0 439.495 0.070 439.845 ;
    RECT 0 439.915 0.070 440.265 ;
    RECT 0 440.335 0.070 440.685 ;
    RECT 0 440.755 0.070 441.105 ;
    RECT 0 441.175 0.070 441.525 ;
    RECT 0 441.595 0.070 441.945 ;
    RECT 0 442.015 0.070 442.365 ;
    RECT 0 442.435 0.070 442.785 ;
    RECT 0 442.855 0.070 443.205 ;
    RECT 0 443.275 0.070 443.625 ;
    RECT 0 443.695 0.070 444.045 ;
    RECT 0 444.115 0.070 444.465 ;
    RECT 0 444.535 0.070 444.885 ;
    RECT 0 444.955 0.070 445.305 ;
    RECT 0 445.375 0.070 445.725 ;
    RECT 0 445.795 0.070 446.145 ;
    RECT 0 446.215 0.070 446.565 ;
    RECT 0 446.635 0.070 446.985 ;
    RECT 0 447.055 0.070 447.405 ;
    RECT 0 447.475 0.070 447.825 ;
    RECT 0 447.895 0.070 448.245 ;
    RECT 0 448.315 0.070 448.665 ;
    RECT 0 448.735 0.070 449.085 ;
    RECT 0 449.155 0.070 449.505 ;
    RECT 0 449.575 0.070 449.925 ;
    RECT 0 449.995 0.070 450.345 ;
    RECT 0 450.415 0.070 450.765 ;
    RECT 0 450.835 0.070 451.185 ;
    RECT 0 451.255 0.070 451.605 ;
    RECT 0 451.675 0.070 452.025 ;
    RECT 0 452.095 0.070 452.445 ;
    RECT 0 452.515 0.070 452.865 ;
    RECT 0 452.935 0.070 453.285 ;
    RECT 0 453.355 0.070 453.705 ;
    RECT 0 453.775 0.070 454.125 ;
    RECT 0 454.195 0.070 454.545 ;
    RECT 0 454.615 0.070 454.965 ;
    RECT 0 455.035 0.070 455.385 ;
    RECT 0 455.455 0.070 455.805 ;
    RECT 0 455.875 0.070 456.225 ;
    RECT 0 456.295 0.070 456.645 ;
    RECT 0 456.715 0.070 457.065 ;
    RECT 0 457.135 0.070 457.485 ;
    RECT 0 457.555 0.070 457.905 ;
    RECT 0 457.975 0.070 458.325 ;
    RECT 0 458.395 0.070 458.745 ;
    RECT 0 458.815 0.070 459.165 ;
    RECT 0 459.235 0.070 487.725 ;
    RECT 0 487.795 0.070 488.145 ;
    RECT 0 488.215 0.070 488.565 ;
    RECT 0 488.635 0.070 488.985 ;
    RECT 0 489.055 0.070 489.405 ;
    RECT 0 489.475 0.070 489.825 ;
    RECT 0 489.895 0.070 490.245 ;
    RECT 0 490.315 0.070 490.665 ;
    RECT 0 490.735 0.070 491.085 ;
    RECT 0 491.155 0.070 491.505 ;
    RECT 0 491.575 0.070 491.925 ;
    RECT 0 491.995 0.070 492.345 ;
    RECT 0 492.415 0.070 492.765 ;
    RECT 0 492.835 0.070 493.185 ;
    RECT 0 493.255 0.070 493.605 ;
    RECT 0 493.675 0.070 494.025 ;
    RECT 0 494.095 0.070 494.445 ;
    RECT 0 494.515 0.070 494.865 ;
    RECT 0 494.935 0.070 495.285 ;
    RECT 0 495.355 0.070 495.705 ;
    RECT 0 495.775 0.070 496.125 ;
    RECT 0 496.195 0.070 496.545 ;
    RECT 0 496.615 0.070 496.965 ;
    RECT 0 497.035 0.070 497.385 ;
    RECT 0 497.455 0.070 497.805 ;
    RECT 0 497.875 0.070 498.225 ;
    RECT 0 498.295 0.070 498.645 ;
    RECT 0 498.715 0.070 499.065 ;
    RECT 0 499.135 0.070 499.485 ;
    RECT 0 499.555 0.070 499.905 ;
    RECT 0 499.975 0.070 500.325 ;
    RECT 0 500.395 0.070 500.745 ;
    RECT 0 500.815 0.070 501.165 ;
    RECT 0 501.235 0.070 501.585 ;
    RECT 0 501.655 0.070 502.005 ;
    RECT 0 502.075 0.070 502.425 ;
    RECT 0 502.495 0.070 502.845 ;
    RECT 0 502.915 0.070 503.265 ;
    RECT 0 503.335 0.070 503.685 ;
    RECT 0 503.755 0.070 504.105 ;
    RECT 0 504.175 0.070 504.525 ;
    RECT 0 504.595 0.070 504.945 ;
    RECT 0 505.015 0.070 505.365 ;
    RECT 0 505.435 0.070 505.785 ;
    RECT 0 505.855 0.070 506.205 ;
    RECT 0 506.275 0.070 506.625 ;
    RECT 0 506.695 0.070 507.045 ;
    RECT 0 507.115 0.070 507.465 ;
    RECT 0 507.535 0.070 507.885 ;
    RECT 0 507.955 0.070 508.305 ;
    RECT 0 508.375 0.070 508.725 ;
    RECT 0 508.795 0.070 509.145 ;
    RECT 0 509.215 0.070 509.565 ;
    RECT 0 509.635 0.070 509.985 ;
    RECT 0 510.055 0.070 510.405 ;
    RECT 0 510.475 0.070 510.825 ;
    RECT 0 510.895 0.070 511.245 ;
    RECT 0 511.315 0.070 511.665 ;
    RECT 0 511.735 0.070 512.085 ;
    RECT 0 512.155 0.070 512.505 ;
    RECT 0 512.575 0.070 512.925 ;
    RECT 0 512.995 0.070 513.345 ;
    RECT 0 513.415 0.070 513.765 ;
    RECT 0 513.835 0.070 514.185 ;
    RECT 0 514.255 0.070 514.605 ;
    RECT 0 514.675 0.070 515.025 ;
    RECT 0 515.095 0.070 515.445 ;
    RECT 0 515.515 0.070 515.865 ;
    RECT 0 515.935 0.070 516.285 ;
    RECT 0 516.355 0.070 516.705 ;
    RECT 0 516.775 0.070 517.125 ;
    RECT 0 517.195 0.070 517.545 ;
    RECT 0 517.615 0.070 517.965 ;
    RECT 0 518.035 0.070 518.385 ;
    RECT 0 518.455 0.070 518.805 ;
    RECT 0 518.875 0.070 519.225 ;
    RECT 0 519.295 0.070 519.645 ;
    RECT 0 519.715 0.070 520.065 ;
    RECT 0 520.135 0.070 520.485 ;
    RECT 0 520.555 0.070 520.905 ;
    RECT 0 520.975 0.070 521.325 ;
    RECT 0 521.395 0.070 521.745 ;
    RECT 0 521.815 0.070 522.165 ;
    RECT 0 522.235 0.070 522.585 ;
    RECT 0 522.655 0.070 523.005 ;
    RECT 0 523.075 0.070 523.425 ;
    RECT 0 523.495 0.070 523.845 ;
    RECT 0 523.915 0.070 524.265 ;
    RECT 0 524.335 0.070 524.685 ;
    RECT 0 524.755 0.070 525.105 ;
    RECT 0 525.175 0.070 525.525 ;
    RECT 0 525.595 0.070 525.945 ;
    RECT 0 526.015 0.070 526.365 ;
    RECT 0 526.435 0.070 526.785 ;
    RECT 0 526.855 0.070 527.205 ;
    RECT 0 527.275 0.070 527.625 ;
    RECT 0 527.695 0.070 528.045 ;
    RECT 0 528.115 0.070 528.465 ;
    RECT 0 528.535 0.070 528.885 ;
    RECT 0 528.955 0.070 529.305 ;
    RECT 0 529.375 0.070 529.725 ;
    RECT 0 529.795 0.070 530.145 ;
    RECT 0 530.215 0.070 530.565 ;
    RECT 0 530.635 0.070 530.985 ;
    RECT 0 531.055 0.070 531.405 ;
    RECT 0 531.475 0.070 531.825 ;
    RECT 0 531.895 0.070 532.245 ;
    RECT 0 532.315 0.070 532.665 ;
    RECT 0 532.735 0.070 533.085 ;
    RECT 0 533.155 0.070 533.505 ;
    RECT 0 533.575 0.070 533.925 ;
    RECT 0 533.995 0.070 534.345 ;
    RECT 0 534.415 0.070 534.765 ;
    RECT 0 534.835 0.070 535.185 ;
    RECT 0 535.255 0.070 535.605 ;
    RECT 0 535.675 0.070 536.025 ;
    RECT 0 536.095 0.070 536.445 ;
    RECT 0 536.515 0.070 536.865 ;
    RECT 0 536.935 0.070 537.285 ;
    RECT 0 537.355 0.070 537.705 ;
    RECT 0 537.775 0.070 538.125 ;
    RECT 0 538.195 0.070 538.545 ;
    RECT 0 538.615 0.070 538.965 ;
    RECT 0 539.035 0.070 539.385 ;
    RECT 0 539.455 0.070 539.805 ;
    RECT 0 539.875 0.070 540.225 ;
    RECT 0 540.295 0.070 540.645 ;
    RECT 0 540.715 0.070 541.065 ;
    RECT 0 541.135 0.070 541.485 ;
    RECT 0 541.555 0.070 541.905 ;
    RECT 0 541.975 0.070 542.325 ;
    RECT 0 542.395 0.070 542.745 ;
    RECT 0 542.815 0.070 543.165 ;
    RECT 0 543.235 0.070 543.585 ;
    RECT 0 543.655 0.070 544.005 ;
    RECT 0 544.075 0.070 544.425 ;
    RECT 0 544.495 0.070 544.845 ;
    RECT 0 544.915 0.070 545.265 ;
    RECT 0 545.335 0.070 545.685 ;
    RECT 0 545.755 0.070 546.105 ;
    RECT 0 546.175 0.070 546.525 ;
    RECT 0 546.595 0.070 546.945 ;
    RECT 0 547.015 0.070 547.365 ;
    RECT 0 547.435 0.070 547.785 ;
    RECT 0 547.855 0.070 548.205 ;
    RECT 0 548.275 0.070 548.625 ;
    RECT 0 548.695 0.070 549.045 ;
    RECT 0 549.115 0.070 549.465 ;
    RECT 0 549.535 0.070 549.885 ;
    RECT 0 549.955 0.070 550.305 ;
    RECT 0 550.375 0.070 550.725 ;
    RECT 0 550.795 0.070 551.145 ;
    RECT 0 551.215 0.070 551.565 ;
    RECT 0 551.635 0.070 551.985 ;
    RECT 0 552.055 0.070 552.405 ;
    RECT 0 552.475 0.070 552.825 ;
    RECT 0 552.895 0.070 553.245 ;
    RECT 0 553.315 0.070 553.665 ;
    RECT 0 553.735 0.070 554.085 ;
    RECT 0 554.155 0.070 554.505 ;
    RECT 0 554.575 0.070 554.925 ;
    RECT 0 554.995 0.070 555.345 ;
    RECT 0 555.415 0.070 555.765 ;
    RECT 0 555.835 0.070 556.185 ;
    RECT 0 556.255 0.070 556.605 ;
    RECT 0 556.675 0.070 557.025 ;
    RECT 0 557.095 0.070 557.445 ;
    RECT 0 557.515 0.070 557.865 ;
    RECT 0 557.935 0.070 558.285 ;
    RECT 0 558.355 0.070 558.705 ;
    RECT 0 558.775 0.070 559.125 ;
    RECT 0 559.195 0.070 559.545 ;
    RECT 0 559.615 0.070 559.965 ;
    RECT 0 560.035 0.070 560.385 ;
    RECT 0 560.455 0.070 560.805 ;
    RECT 0 560.875 0.070 561.225 ;
    RECT 0 561.295 0.070 561.645 ;
    RECT 0 561.715 0.070 562.065 ;
    RECT 0 562.135 0.070 562.485 ;
    RECT 0 562.555 0.070 562.905 ;
    RECT 0 562.975 0.070 563.325 ;
    RECT 0 563.395 0.070 563.745 ;
    RECT 0 563.815 0.070 564.165 ;
    RECT 0 564.235 0.070 564.585 ;
    RECT 0 564.655 0.070 565.005 ;
    RECT 0 565.075 0.070 565.425 ;
    RECT 0 565.495 0.070 565.845 ;
    RECT 0 565.915 0.070 566.265 ;
    RECT 0 566.335 0.070 566.685 ;
    RECT 0 566.755 0.070 567.105 ;
    RECT 0 567.175 0.070 567.525 ;
    RECT 0 567.595 0.070 567.945 ;
    RECT 0 568.015 0.070 568.365 ;
    RECT 0 568.435 0.070 568.785 ;
    RECT 0 568.855 0.070 569.205 ;
    RECT 0 569.275 0.070 569.625 ;
    RECT 0 569.695 0.070 570.045 ;
    RECT 0 570.115 0.070 570.465 ;
    RECT 0 570.535 0.070 570.885 ;
    RECT 0 570.955 0.070 571.305 ;
    RECT 0 571.375 0.070 571.725 ;
    RECT 0 571.795 0.070 572.145 ;
    RECT 0 572.215 0.070 572.565 ;
    RECT 0 572.635 0.070 572.985 ;
    RECT 0 573.055 0.070 573.405 ;
    RECT 0 573.475 0.070 573.825 ;
    RECT 0 573.895 0.070 574.245 ;
    RECT 0 574.315 0.070 574.665 ;
    RECT 0 574.735 0.070 575.085 ;
    RECT 0 575.155 0.070 575.505 ;
    RECT 0 575.575 0.070 575.925 ;
    RECT 0 575.995 0.070 576.345 ;
    RECT 0 576.415 0.070 576.765 ;
    RECT 0 576.835 0.070 577.185 ;
    RECT 0 577.255 0.070 577.605 ;
    RECT 0 577.675 0.070 578.025 ;
    RECT 0 578.095 0.070 578.445 ;
    RECT 0 578.515 0.070 578.865 ;
    RECT 0 578.935 0.070 579.285 ;
    RECT 0 579.355 0.070 579.705 ;
    RECT 0 579.775 0.070 580.125 ;
    RECT 0 580.195 0.070 580.545 ;
    RECT 0 580.615 0.070 580.965 ;
    RECT 0 581.035 0.070 581.385 ;
    RECT 0 581.455 0.070 581.805 ;
    RECT 0 581.875 0.070 582.225 ;
    RECT 0 582.295 0.070 582.645 ;
    RECT 0 582.715 0.070 583.065 ;
    RECT 0 583.135 0.070 583.485 ;
    RECT 0 583.555 0.070 583.905 ;
    RECT 0 583.975 0.070 584.325 ;
    RECT 0 584.395 0.070 584.745 ;
    RECT 0 584.815 0.070 585.165 ;
    RECT 0 585.235 0.070 585.585 ;
    RECT 0 585.655 0.070 586.005 ;
    RECT 0 586.075 0.070 586.425 ;
    RECT 0 586.495 0.070 586.845 ;
    RECT 0 586.915 0.070 587.265 ;
    RECT 0 587.335 0.070 587.685 ;
    RECT 0 587.755 0.070 588.105 ;
    RECT 0 588.175 0.070 588.525 ;
    RECT 0 588.595 0.070 588.945 ;
    RECT 0 589.015 0.070 589.365 ;
    RECT 0 589.435 0.070 589.785 ;
    RECT 0 589.855 0.070 590.205 ;
    RECT 0 590.275 0.070 590.625 ;
    RECT 0 590.695 0.070 591.045 ;
    RECT 0 591.115 0.070 591.465 ;
    RECT 0 591.535 0.070 591.885 ;
    RECT 0 591.955 0.070 592.305 ;
    RECT 0 592.375 0.070 592.725 ;
    RECT 0 592.795 0.070 593.145 ;
    RECT 0 593.215 0.070 593.565 ;
    RECT 0 593.635 0.070 593.985 ;
    RECT 0 594.055 0.070 594.405 ;
    RECT 0 594.475 0.070 594.825 ;
    RECT 0 594.895 0.070 595.245 ;
    RECT 0 595.315 0.070 595.665 ;
    RECT 0 595.735 0.070 596.085 ;
    RECT 0 596.155 0.070 596.505 ;
    RECT 0 596.575 0.070 596.925 ;
    RECT 0 596.995 0.070 597.345 ;
    RECT 0 597.415 0.070 597.765 ;
    RECT 0 597.835 0.070 598.185 ;
    RECT 0 598.255 0.070 598.605 ;
    RECT 0 598.675 0.070 599.025 ;
    RECT 0 599.095 0.070 599.445 ;
    RECT 0 599.515 0.070 599.865 ;
    RECT 0 599.935 0.070 600.285 ;
    RECT 0 600.355 0.070 600.705 ;
    RECT 0 600.775 0.070 601.125 ;
    RECT 0 601.195 0.070 601.545 ;
    RECT 0 601.615 0.070 601.965 ;
    RECT 0 602.035 0.070 602.385 ;
    RECT 0 602.455 0.070 602.805 ;
    RECT 0 602.875 0.070 603.225 ;
    RECT 0 603.295 0.070 603.645 ;
    RECT 0 603.715 0.070 604.065 ;
    RECT 0 604.135 0.070 604.485 ;
    RECT 0 604.555 0.070 604.905 ;
    RECT 0 604.975 0.070 605.325 ;
    RECT 0 605.395 0.070 605.745 ;
    RECT 0 605.815 0.070 606.165 ;
    RECT 0 606.235 0.070 606.585 ;
    RECT 0 606.655 0.070 607.005 ;
    RECT 0 607.075 0.070 607.425 ;
    RECT 0 607.495 0.070 607.845 ;
    RECT 0 607.915 0.070 608.265 ;
    RECT 0 608.335 0.070 608.685 ;
    RECT 0 608.755 0.070 609.105 ;
    RECT 0 609.175 0.070 609.525 ;
    RECT 0 609.595 0.070 609.945 ;
    RECT 0 610.015 0.070 610.365 ;
    RECT 0 610.435 0.070 610.785 ;
    RECT 0 610.855 0.070 611.205 ;
    RECT 0 611.275 0.070 611.625 ;
    RECT 0 611.695 0.070 612.045 ;
    RECT 0 612.115 0.070 612.465 ;
    RECT 0 612.535 0.070 612.885 ;
    RECT 0 612.955 0.070 613.305 ;
    RECT 0 613.375 0.070 613.725 ;
    RECT 0 613.795 0.070 614.145 ;
    RECT 0 614.215 0.070 614.565 ;
    RECT 0 614.635 0.070 614.985 ;
    RECT 0 615.055 0.070 615.405 ;
    RECT 0 615.475 0.070 615.825 ;
    RECT 0 615.895 0.070 616.245 ;
    RECT 0 616.315 0.070 616.665 ;
    RECT 0 616.735 0.070 617.085 ;
    RECT 0 617.155 0.070 617.505 ;
    RECT 0 617.575 0.070 617.925 ;
    RECT 0 617.995 0.070 618.345 ;
    RECT 0 618.415 0.070 618.765 ;
    RECT 0 618.835 0.070 619.185 ;
    RECT 0 619.255 0.070 619.605 ;
    RECT 0 619.675 0.070 620.025 ;
    RECT 0 620.095 0.070 620.445 ;
    RECT 0 620.515 0.070 620.865 ;
    RECT 0 620.935 0.070 621.285 ;
    RECT 0 621.355 0.070 621.705 ;
    RECT 0 621.775 0.070 622.125 ;
    RECT 0 622.195 0.070 622.545 ;
    RECT 0 622.615 0.070 622.965 ;
    RECT 0 623.035 0.070 623.385 ;
    RECT 0 623.455 0.070 623.805 ;
    RECT 0 623.875 0.070 624.225 ;
    RECT 0 624.295 0.070 624.645 ;
    RECT 0 624.715 0.070 625.065 ;
    RECT 0 625.135 0.070 625.485 ;
    RECT 0 625.555 0.070 625.905 ;
    RECT 0 625.975 0.070 626.325 ;
    RECT 0 626.395 0.070 626.745 ;
    RECT 0 626.815 0.070 627.165 ;
    RECT 0 627.235 0.070 627.585 ;
    RECT 0 627.655 0.070 628.005 ;
    RECT 0 628.075 0.070 628.425 ;
    RECT 0 628.495 0.070 628.845 ;
    RECT 0 628.915 0.070 629.265 ;
    RECT 0 629.335 0.070 629.685 ;
    RECT 0 629.755 0.070 630.105 ;
    RECT 0 630.175 0.070 630.525 ;
    RECT 0 630.595 0.070 630.945 ;
    RECT 0 631.015 0.070 631.365 ;
    RECT 0 631.435 0.070 631.785 ;
    RECT 0 631.855 0.070 632.205 ;
    RECT 0 632.275 0.070 632.625 ;
    RECT 0 632.695 0.070 633.045 ;
    RECT 0 633.115 0.070 633.465 ;
    RECT 0 633.535 0.070 633.885 ;
    RECT 0 633.955 0.070 634.305 ;
    RECT 0 634.375 0.070 634.725 ;
    RECT 0 634.795 0.070 635.145 ;
    RECT 0 635.215 0.070 635.565 ;
    RECT 0 635.635 0.070 635.985 ;
    RECT 0 636.055 0.070 636.405 ;
    RECT 0 636.475 0.070 636.825 ;
    RECT 0 636.895 0.070 637.245 ;
    RECT 0 637.315 0.070 637.665 ;
    RECT 0 637.735 0.070 638.085 ;
    RECT 0 638.155 0.070 638.505 ;
    RECT 0 638.575 0.070 638.925 ;
    RECT 0 638.995 0.070 639.345 ;
    RECT 0 639.415 0.070 639.765 ;
    RECT 0 639.835 0.070 640.185 ;
    RECT 0 640.255 0.070 640.605 ;
    RECT 0 640.675 0.070 641.025 ;
    RECT 0 641.095 0.070 641.445 ;
    RECT 0 641.515 0.070 641.865 ;
    RECT 0 641.935 0.070 642.285 ;
    RECT 0 642.355 0.070 642.705 ;
    RECT 0 642.775 0.070 643.125 ;
    RECT 0 643.195 0.070 643.545 ;
    RECT 0 643.615 0.070 643.965 ;
    RECT 0 644.035 0.070 644.385 ;
    RECT 0 644.455 0.070 644.805 ;
    RECT 0 644.875 0.070 645.225 ;
    RECT 0 645.295 0.070 645.645 ;
    RECT 0 645.715 0.070 646.065 ;
    RECT 0 646.135 0.070 646.485 ;
    RECT 0 646.555 0.070 646.905 ;
    RECT 0 646.975 0.070 647.325 ;
    RECT 0 647.395 0.070 647.745 ;
    RECT 0 647.815 0.070 648.165 ;
    RECT 0 648.235 0.070 648.585 ;
    RECT 0 648.655 0.070 649.005 ;
    RECT 0 649.075 0.070 649.425 ;
    RECT 0 649.495 0.070 649.845 ;
    RECT 0 649.915 0.070 650.265 ;
    RECT 0 650.335 0.070 650.685 ;
    RECT 0 650.755 0.070 651.105 ;
    RECT 0 651.175 0.070 651.525 ;
    RECT 0 651.595 0.070 651.945 ;
    RECT 0 652.015 0.070 652.365 ;
    RECT 0 652.435 0.070 652.785 ;
    RECT 0 652.855 0.070 653.205 ;
    RECT 0 653.275 0.070 653.625 ;
    RECT 0 653.695 0.070 654.045 ;
    RECT 0 654.115 0.070 654.465 ;
    RECT 0 654.535 0.070 654.885 ;
    RECT 0 654.955 0.070 655.305 ;
    RECT 0 655.375 0.070 655.725 ;
    RECT 0 655.795 0.070 656.145 ;
    RECT 0 656.215 0.070 656.565 ;
    RECT 0 656.635 0.070 656.985 ;
    RECT 0 657.055 0.070 657.405 ;
    RECT 0 657.475 0.070 657.825 ;
    RECT 0 657.895 0.070 658.245 ;
    RECT 0 658.315 0.070 658.665 ;
    RECT 0 658.735 0.070 659.085 ;
    RECT 0 659.155 0.070 659.505 ;
    RECT 0 659.575 0.070 659.925 ;
    RECT 0 659.995 0.070 660.345 ;
    RECT 0 660.415 0.070 660.765 ;
    RECT 0 660.835 0.070 661.185 ;
    RECT 0 661.255 0.070 661.605 ;
    RECT 0 661.675 0.070 662.025 ;
    RECT 0 662.095 0.070 662.445 ;
    RECT 0 662.515 0.070 662.865 ;
    RECT 0 662.935 0.070 663.285 ;
    RECT 0 663.355 0.070 663.705 ;
    RECT 0 663.775 0.070 664.125 ;
    RECT 0 664.195 0.070 664.545 ;
    RECT 0 664.615 0.070 664.965 ;
    RECT 0 665.035 0.070 665.385 ;
    RECT 0 665.455 0.070 665.805 ;
    RECT 0 665.875 0.070 666.225 ;
    RECT 0 666.295 0.070 666.645 ;
    RECT 0 666.715 0.070 667.065 ;
    RECT 0 667.135 0.070 667.485 ;
    RECT 0 667.555 0.070 667.905 ;
    RECT 0 667.975 0.070 668.325 ;
    RECT 0 668.395 0.070 668.745 ;
    RECT 0 668.815 0.070 669.165 ;
    RECT 0 669.235 0.070 669.585 ;
    RECT 0 669.655 0.070 670.005 ;
    RECT 0 670.075 0.070 670.425 ;
    RECT 0 670.495 0.070 670.845 ;
    RECT 0 670.915 0.070 671.265 ;
    RECT 0 671.335 0.070 671.685 ;
    RECT 0 671.755 0.070 672.105 ;
    RECT 0 672.175 0.070 672.525 ;
    RECT 0 672.595 0.070 672.945 ;
    RECT 0 673.015 0.070 673.365 ;
    RECT 0 673.435 0.070 673.785 ;
    RECT 0 673.855 0.070 674.205 ;
    RECT 0 674.275 0.070 674.625 ;
    RECT 0 674.695 0.070 675.045 ;
    RECT 0 675.115 0.070 675.465 ;
    RECT 0 675.535 0.070 675.885 ;
    RECT 0 675.955 0.070 676.305 ;
    RECT 0 676.375 0.070 676.725 ;
    RECT 0 676.795 0.070 677.145 ;
    RECT 0 677.215 0.070 677.565 ;
    RECT 0 677.635 0.070 677.985 ;
    RECT 0 678.055 0.070 678.405 ;
    RECT 0 678.475 0.070 678.825 ;
    RECT 0 678.895 0.070 679.245 ;
    RECT 0 679.315 0.070 679.665 ;
    RECT 0 679.735 0.070 680.085 ;
    RECT 0 680.155 0.070 680.505 ;
    RECT 0 680.575 0.070 680.925 ;
    RECT 0 680.995 0.070 681.345 ;
    RECT 0 681.415 0.070 681.765 ;
    RECT 0 681.835 0.070 682.185 ;
    RECT 0 682.255 0.070 682.605 ;
    RECT 0 682.675 0.070 683.025 ;
    RECT 0 683.095 0.070 683.445 ;
    RECT 0 683.515 0.070 683.865 ;
    RECT 0 683.935 0.070 684.285 ;
    RECT 0 684.355 0.070 684.705 ;
    RECT 0 684.775 0.070 685.125 ;
    RECT 0 685.195 0.070 685.545 ;
    RECT 0 685.615 0.070 685.965 ;
    RECT 0 686.035 0.070 686.385 ;
    RECT 0 686.455 0.070 686.805 ;
    RECT 0 686.875 0.070 687.225 ;
    RECT 0 687.295 0.070 687.645 ;
    RECT 0 687.715 0.070 688.065 ;
    RECT 0 688.135 0.070 688.485 ;
    RECT 0 688.555 0.070 688.905 ;
    RECT 0 688.975 0.070 689.325 ;
    RECT 0 689.395 0.070 689.745 ;
    RECT 0 689.815 0.070 690.165 ;
    RECT 0 690.235 0.070 690.585 ;
    RECT 0 690.655 0.070 691.005 ;
    RECT 0 691.075 0.070 691.425 ;
    RECT 0 691.495 0.070 691.845 ;
    RECT 0 691.915 0.070 692.265 ;
    RECT 0 692.335 0.070 692.685 ;
    RECT 0 692.755 0.070 693.105 ;
    RECT 0 693.175 0.070 693.525 ;
    RECT 0 693.595 0.070 693.945 ;
    RECT 0 694.015 0.070 694.365 ;
    RECT 0 694.435 0.070 694.785 ;
    RECT 0 694.855 0.070 695.205 ;
    RECT 0 695.275 0.070 695.625 ;
    RECT 0 695.695 0.070 696.045 ;
    RECT 0 696.115 0.070 696.465 ;
    RECT 0 696.535 0.070 696.885 ;
    RECT 0 696.955 0.070 697.305 ;
    RECT 0 697.375 0.070 697.725 ;
    RECT 0 697.795 0.070 698.145 ;
    RECT 0 698.215 0.070 698.565 ;
    RECT 0 698.635 0.070 698.985 ;
    RECT 0 699.055 0.070 699.405 ;
    RECT 0 699.475 0.070 699.825 ;
    RECT 0 699.895 0.070 700.245 ;
    RECT 0 700.315 0.070 700.665 ;
    RECT 0 700.735 0.070 701.085 ;
    RECT 0 701.155 0.070 701.505 ;
    RECT 0 701.575 0.070 701.925 ;
    RECT 0 701.995 0.070 702.345 ;
    RECT 0 702.415 0.070 730.905 ;
    RECT 0 730.975 0.070 731.325 ;
    RECT 0 731.395 0.070 731.745 ;
    RECT 0 731.815 0.070 732.165 ;
    RECT 0 732.235 0.070 732.585 ;
    RECT 0 732.655 0.070 733.005 ;
    RECT 0 733.075 0.070 733.425 ;
    RECT 0 733.495 0.070 733.845 ;
    RECT 0 733.915 0.070 762.405 ;
    RECT 0 762.475 0.070 762.825 ;
    RECT 0 762.895 0.070 763.245 ;
    RECT 0 763.315 0.070 767.200 ;
    LAYER metal4 ;
    RECT 0 0 689.130 1.400 ;
    RECT 0 765.800 689.130 767.200 ;
    RECT 0.000 1.400 1.260 765.800 ;
    RECT 1.540 1.400 2.380 765.800 ;
    RECT 2.660 1.400 3.500 765.800 ;
    RECT 3.780 1.400 4.620 765.800 ;
    RECT 4.900 1.400 5.740 765.800 ;
    RECT 6.020 1.400 6.860 765.800 ;
    RECT 7.140 1.400 7.980 765.800 ;
    RECT 8.260 1.400 9.100 765.800 ;
    RECT 9.380 1.400 10.220 765.800 ;
    RECT 10.500 1.400 11.340 765.800 ;
    RECT 11.620 1.400 12.460 765.800 ;
    RECT 12.740 1.400 13.580 765.800 ;
    RECT 13.860 1.400 14.700 765.800 ;
    RECT 14.980 1.400 15.820 765.800 ;
    RECT 16.100 1.400 16.940 765.800 ;
    RECT 17.220 1.400 18.060 765.800 ;
    RECT 18.340 1.400 19.180 765.800 ;
    RECT 19.460 1.400 20.300 765.800 ;
    RECT 20.580 1.400 21.420 765.800 ;
    RECT 21.700 1.400 22.540 765.800 ;
    RECT 22.820 1.400 23.660 765.800 ;
    RECT 23.940 1.400 24.780 765.800 ;
    RECT 25.060 1.400 25.900 765.800 ;
    RECT 26.180 1.400 27.020 765.800 ;
    RECT 27.300 1.400 28.140 765.800 ;
    RECT 28.420 1.400 29.260 765.800 ;
    RECT 29.540 1.400 30.380 765.800 ;
    RECT 30.660 1.400 31.500 765.800 ;
    RECT 31.780 1.400 32.620 765.800 ;
    RECT 32.900 1.400 33.740 765.800 ;
    RECT 34.020 1.400 34.860 765.800 ;
    RECT 35.140 1.400 35.980 765.800 ;
    RECT 36.260 1.400 37.100 765.800 ;
    RECT 37.380 1.400 38.220 765.800 ;
    RECT 38.500 1.400 39.340 765.800 ;
    RECT 39.620 1.400 40.460 765.800 ;
    RECT 40.740 1.400 41.580 765.800 ;
    RECT 41.860 1.400 42.700 765.800 ;
    RECT 42.980 1.400 43.820 765.800 ;
    RECT 44.100 1.400 44.940 765.800 ;
    RECT 45.220 1.400 46.060 765.800 ;
    RECT 46.340 1.400 47.180 765.800 ;
    RECT 47.460 1.400 48.300 765.800 ;
    RECT 48.580 1.400 49.420 765.800 ;
    RECT 49.700 1.400 50.540 765.800 ;
    RECT 50.820 1.400 51.660 765.800 ;
    RECT 51.940 1.400 52.780 765.800 ;
    RECT 53.060 1.400 53.900 765.800 ;
    RECT 54.180 1.400 55.020 765.800 ;
    RECT 55.300 1.400 56.140 765.800 ;
    RECT 56.420 1.400 57.260 765.800 ;
    RECT 57.540 1.400 58.380 765.800 ;
    RECT 58.660 1.400 59.500 765.800 ;
    RECT 59.780 1.400 60.620 765.800 ;
    RECT 60.900 1.400 61.740 765.800 ;
    RECT 62.020 1.400 62.860 765.800 ;
    RECT 63.140 1.400 63.980 765.800 ;
    RECT 64.260 1.400 65.100 765.800 ;
    RECT 65.380 1.400 66.220 765.800 ;
    RECT 66.500 1.400 67.340 765.800 ;
    RECT 67.620 1.400 68.460 765.800 ;
    RECT 68.740 1.400 69.580 765.800 ;
    RECT 69.860 1.400 70.700 765.800 ;
    RECT 70.980 1.400 71.820 765.800 ;
    RECT 72.100 1.400 72.940 765.800 ;
    RECT 73.220 1.400 74.060 765.800 ;
    RECT 74.340 1.400 75.180 765.800 ;
    RECT 75.460 1.400 76.300 765.800 ;
    RECT 76.580 1.400 77.420 765.800 ;
    RECT 77.700 1.400 78.540 765.800 ;
    RECT 78.820 1.400 79.660 765.800 ;
    RECT 79.940 1.400 80.780 765.800 ;
    RECT 81.060 1.400 81.900 765.800 ;
    RECT 82.180 1.400 83.020 765.800 ;
    RECT 83.300 1.400 84.140 765.800 ;
    RECT 84.420 1.400 85.260 765.800 ;
    RECT 85.540 1.400 86.380 765.800 ;
    RECT 86.660 1.400 87.500 765.800 ;
    RECT 87.780 1.400 88.620 765.800 ;
    RECT 88.900 1.400 89.740 765.800 ;
    RECT 90.020 1.400 90.860 765.800 ;
    RECT 91.140 1.400 91.980 765.800 ;
    RECT 92.260 1.400 93.100 765.800 ;
    RECT 93.380 1.400 94.220 765.800 ;
    RECT 94.500 1.400 95.340 765.800 ;
    RECT 95.620 1.400 96.460 765.800 ;
    RECT 96.740 1.400 97.580 765.800 ;
    RECT 97.860 1.400 98.700 765.800 ;
    RECT 98.980 1.400 99.820 765.800 ;
    RECT 100.100 1.400 100.940 765.800 ;
    RECT 101.220 1.400 102.060 765.800 ;
    RECT 102.340 1.400 103.180 765.800 ;
    RECT 103.460 1.400 104.300 765.800 ;
    RECT 104.580 1.400 105.420 765.800 ;
    RECT 105.700 1.400 106.540 765.800 ;
    RECT 106.820 1.400 107.660 765.800 ;
    RECT 107.940 1.400 108.780 765.800 ;
    RECT 109.060 1.400 109.900 765.800 ;
    RECT 110.180 1.400 111.020 765.800 ;
    RECT 111.300 1.400 112.140 765.800 ;
    RECT 112.420 1.400 113.260 765.800 ;
    RECT 113.540 1.400 114.380 765.800 ;
    RECT 114.660 1.400 115.500 765.800 ;
    RECT 115.780 1.400 116.620 765.800 ;
    RECT 116.900 1.400 117.740 765.800 ;
    RECT 118.020 1.400 118.860 765.800 ;
    RECT 119.140 1.400 119.980 765.800 ;
    RECT 120.260 1.400 121.100 765.800 ;
    RECT 121.380 1.400 122.220 765.800 ;
    RECT 122.500 1.400 123.340 765.800 ;
    RECT 123.620 1.400 124.460 765.800 ;
    RECT 124.740 1.400 125.580 765.800 ;
    RECT 125.860 1.400 126.700 765.800 ;
    RECT 126.980 1.400 127.820 765.800 ;
    RECT 128.100 1.400 128.940 765.800 ;
    RECT 129.220 1.400 130.060 765.800 ;
    RECT 130.340 1.400 131.180 765.800 ;
    RECT 131.460 1.400 132.300 765.800 ;
    RECT 132.580 1.400 133.420 765.800 ;
    RECT 133.700 1.400 134.540 765.800 ;
    RECT 134.820 1.400 135.660 765.800 ;
    RECT 135.940 1.400 136.780 765.800 ;
    RECT 137.060 1.400 137.900 765.800 ;
    RECT 138.180 1.400 139.020 765.800 ;
    RECT 139.300 1.400 140.140 765.800 ;
    RECT 140.420 1.400 141.260 765.800 ;
    RECT 141.540 1.400 142.380 765.800 ;
    RECT 142.660 1.400 143.500 765.800 ;
    RECT 143.780 1.400 144.620 765.800 ;
    RECT 144.900 1.400 145.740 765.800 ;
    RECT 146.020 1.400 146.860 765.800 ;
    RECT 147.140 1.400 147.980 765.800 ;
    RECT 148.260 1.400 149.100 765.800 ;
    RECT 149.380 1.400 150.220 765.800 ;
    RECT 150.500 1.400 151.340 765.800 ;
    RECT 151.620 1.400 152.460 765.800 ;
    RECT 152.740 1.400 153.580 765.800 ;
    RECT 153.860 1.400 154.700 765.800 ;
    RECT 154.980 1.400 155.820 765.800 ;
    RECT 156.100 1.400 156.940 765.800 ;
    RECT 157.220 1.400 158.060 765.800 ;
    RECT 158.340 1.400 159.180 765.800 ;
    RECT 159.460 1.400 160.300 765.800 ;
    RECT 160.580 1.400 161.420 765.800 ;
    RECT 161.700 1.400 162.540 765.800 ;
    RECT 162.820 1.400 163.660 765.800 ;
    RECT 163.940 1.400 164.780 765.800 ;
    RECT 165.060 1.400 165.900 765.800 ;
    RECT 166.180 1.400 167.020 765.800 ;
    RECT 167.300 1.400 168.140 765.800 ;
    RECT 168.420 1.400 169.260 765.800 ;
    RECT 169.540 1.400 170.380 765.800 ;
    RECT 170.660 1.400 171.500 765.800 ;
    RECT 171.780 1.400 172.620 765.800 ;
    RECT 172.900 1.400 173.740 765.800 ;
    RECT 174.020 1.400 174.860 765.800 ;
    RECT 175.140 1.400 175.980 765.800 ;
    RECT 176.260 1.400 177.100 765.800 ;
    RECT 177.380 1.400 178.220 765.800 ;
    RECT 178.500 1.400 179.340 765.800 ;
    RECT 179.620 1.400 180.460 765.800 ;
    RECT 180.740 1.400 181.580 765.800 ;
    RECT 181.860 1.400 182.700 765.800 ;
    RECT 182.980 1.400 183.820 765.800 ;
    RECT 184.100 1.400 184.940 765.800 ;
    RECT 185.220 1.400 186.060 765.800 ;
    RECT 186.340 1.400 187.180 765.800 ;
    RECT 187.460 1.400 188.300 765.800 ;
    RECT 188.580 1.400 189.420 765.800 ;
    RECT 189.700 1.400 190.540 765.800 ;
    RECT 190.820 1.400 191.660 765.800 ;
    RECT 191.940 1.400 192.780 765.800 ;
    RECT 193.060 1.400 193.900 765.800 ;
    RECT 194.180 1.400 195.020 765.800 ;
    RECT 195.300 1.400 196.140 765.800 ;
    RECT 196.420 1.400 197.260 765.800 ;
    RECT 197.540 1.400 198.380 765.800 ;
    RECT 198.660 1.400 199.500 765.800 ;
    RECT 199.780 1.400 200.620 765.800 ;
    RECT 200.900 1.400 201.740 765.800 ;
    RECT 202.020 1.400 202.860 765.800 ;
    RECT 203.140 1.400 203.980 765.800 ;
    RECT 204.260 1.400 205.100 765.800 ;
    RECT 205.380 1.400 206.220 765.800 ;
    RECT 206.500 1.400 207.340 765.800 ;
    RECT 207.620 1.400 208.460 765.800 ;
    RECT 208.740 1.400 209.580 765.800 ;
    RECT 209.860 1.400 210.700 765.800 ;
    RECT 210.980 1.400 211.820 765.800 ;
    RECT 212.100 1.400 212.940 765.800 ;
    RECT 213.220 1.400 214.060 765.800 ;
    RECT 214.340 1.400 215.180 765.800 ;
    RECT 215.460 1.400 216.300 765.800 ;
    RECT 216.580 1.400 217.420 765.800 ;
    RECT 217.700 1.400 218.540 765.800 ;
    RECT 218.820 1.400 219.660 765.800 ;
    RECT 219.940 1.400 220.780 765.800 ;
    RECT 221.060 1.400 221.900 765.800 ;
    RECT 222.180 1.400 223.020 765.800 ;
    RECT 223.300 1.400 224.140 765.800 ;
    RECT 224.420 1.400 225.260 765.800 ;
    RECT 225.540 1.400 226.380 765.800 ;
    RECT 226.660 1.400 227.500 765.800 ;
    RECT 227.780 1.400 228.620 765.800 ;
    RECT 228.900 1.400 229.740 765.800 ;
    RECT 230.020 1.400 230.860 765.800 ;
    RECT 231.140 1.400 231.980 765.800 ;
    RECT 232.260 1.400 233.100 765.800 ;
    RECT 233.380 1.400 234.220 765.800 ;
    RECT 234.500 1.400 235.340 765.800 ;
    RECT 235.620 1.400 236.460 765.800 ;
    RECT 236.740 1.400 237.580 765.800 ;
    RECT 237.860 1.400 238.700 765.800 ;
    RECT 238.980 1.400 239.820 765.800 ;
    RECT 240.100 1.400 240.940 765.800 ;
    RECT 241.220 1.400 242.060 765.800 ;
    RECT 242.340 1.400 243.180 765.800 ;
    RECT 243.460 1.400 244.300 765.800 ;
    RECT 244.580 1.400 245.420 765.800 ;
    RECT 245.700 1.400 246.540 765.800 ;
    RECT 246.820 1.400 247.660 765.800 ;
    RECT 247.940 1.400 248.780 765.800 ;
    RECT 249.060 1.400 249.900 765.800 ;
    RECT 250.180 1.400 251.020 765.800 ;
    RECT 251.300 1.400 252.140 765.800 ;
    RECT 252.420 1.400 253.260 765.800 ;
    RECT 253.540 1.400 254.380 765.800 ;
    RECT 254.660 1.400 255.500 765.800 ;
    RECT 255.780 1.400 256.620 765.800 ;
    RECT 256.900 1.400 257.740 765.800 ;
    RECT 258.020 1.400 258.860 765.800 ;
    RECT 259.140 1.400 259.980 765.800 ;
    RECT 260.260 1.400 261.100 765.800 ;
    RECT 261.380 1.400 262.220 765.800 ;
    RECT 262.500 1.400 263.340 765.800 ;
    RECT 263.620 1.400 264.460 765.800 ;
    RECT 264.740 1.400 265.580 765.800 ;
    RECT 265.860 1.400 266.700 765.800 ;
    RECT 266.980 1.400 267.820 765.800 ;
    RECT 268.100 1.400 268.940 765.800 ;
    RECT 269.220 1.400 270.060 765.800 ;
    RECT 270.340 1.400 271.180 765.800 ;
    RECT 271.460 1.400 272.300 765.800 ;
    RECT 272.580 1.400 273.420 765.800 ;
    RECT 273.700 1.400 274.540 765.800 ;
    RECT 274.820 1.400 275.660 765.800 ;
    RECT 275.940 1.400 276.780 765.800 ;
    RECT 277.060 1.400 277.900 765.800 ;
    RECT 278.180 1.400 279.020 765.800 ;
    RECT 279.300 1.400 280.140 765.800 ;
    RECT 280.420 1.400 281.260 765.800 ;
    RECT 281.540 1.400 282.380 765.800 ;
    RECT 282.660 1.400 283.500 765.800 ;
    RECT 283.780 1.400 284.620 765.800 ;
    RECT 284.900 1.400 285.740 765.800 ;
    RECT 286.020 1.400 286.860 765.800 ;
    RECT 287.140 1.400 287.980 765.800 ;
    RECT 288.260 1.400 289.100 765.800 ;
    RECT 289.380 1.400 290.220 765.800 ;
    RECT 290.500 1.400 291.340 765.800 ;
    RECT 291.620 1.400 292.460 765.800 ;
    RECT 292.740 1.400 293.580 765.800 ;
    RECT 293.860 1.400 294.700 765.800 ;
    RECT 294.980 1.400 295.820 765.800 ;
    RECT 296.100 1.400 296.940 765.800 ;
    RECT 297.220 1.400 298.060 765.800 ;
    RECT 298.340 1.400 299.180 765.800 ;
    RECT 299.460 1.400 300.300 765.800 ;
    RECT 300.580 1.400 301.420 765.800 ;
    RECT 301.700 1.400 302.540 765.800 ;
    RECT 302.820 1.400 303.660 765.800 ;
    RECT 303.940 1.400 304.780 765.800 ;
    RECT 305.060 1.400 305.900 765.800 ;
    RECT 306.180 1.400 307.020 765.800 ;
    RECT 307.300 1.400 308.140 765.800 ;
    RECT 308.420 1.400 309.260 765.800 ;
    RECT 309.540 1.400 310.380 765.800 ;
    RECT 310.660 1.400 311.500 765.800 ;
    RECT 311.780 1.400 312.620 765.800 ;
    RECT 312.900 1.400 313.740 765.800 ;
    RECT 314.020 1.400 314.860 765.800 ;
    RECT 315.140 1.400 315.980 765.800 ;
    RECT 316.260 1.400 317.100 765.800 ;
    RECT 317.380 1.400 318.220 765.800 ;
    RECT 318.500 1.400 319.340 765.800 ;
    RECT 319.620 1.400 320.460 765.800 ;
    RECT 320.740 1.400 321.580 765.800 ;
    RECT 321.860 1.400 322.700 765.800 ;
    RECT 322.980 1.400 323.820 765.800 ;
    RECT 324.100 1.400 324.940 765.800 ;
    RECT 325.220 1.400 326.060 765.800 ;
    RECT 326.340 1.400 327.180 765.800 ;
    RECT 327.460 1.400 328.300 765.800 ;
    RECT 328.580 1.400 329.420 765.800 ;
    RECT 329.700 1.400 330.540 765.800 ;
    RECT 330.820 1.400 331.660 765.800 ;
    RECT 331.940 1.400 332.780 765.800 ;
    RECT 333.060 1.400 333.900 765.800 ;
    RECT 334.180 1.400 335.020 765.800 ;
    RECT 335.300 1.400 336.140 765.800 ;
    RECT 336.420 1.400 337.260 765.800 ;
    RECT 337.540 1.400 338.380 765.800 ;
    RECT 338.660 1.400 339.500 765.800 ;
    RECT 339.780 1.400 340.620 765.800 ;
    RECT 340.900 1.400 341.740 765.800 ;
    RECT 342.020 1.400 342.860 765.800 ;
    RECT 343.140 1.400 343.980 765.800 ;
    RECT 344.260 1.400 345.100 765.800 ;
    RECT 345.380 1.400 346.220 765.800 ;
    RECT 346.500 1.400 347.340 765.800 ;
    RECT 347.620 1.400 348.460 765.800 ;
    RECT 348.740 1.400 349.580 765.800 ;
    RECT 349.860 1.400 350.700 765.800 ;
    RECT 350.980 1.400 351.820 765.800 ;
    RECT 352.100 1.400 352.940 765.800 ;
    RECT 353.220 1.400 354.060 765.800 ;
    RECT 354.340 1.400 355.180 765.800 ;
    RECT 355.460 1.400 356.300 765.800 ;
    RECT 356.580 1.400 357.420 765.800 ;
    RECT 357.700 1.400 358.540 765.800 ;
    RECT 358.820 1.400 359.660 765.800 ;
    RECT 359.940 1.400 360.780 765.800 ;
    RECT 361.060 1.400 361.900 765.800 ;
    RECT 362.180 1.400 363.020 765.800 ;
    RECT 363.300 1.400 364.140 765.800 ;
    RECT 364.420 1.400 365.260 765.800 ;
    RECT 365.540 1.400 366.380 765.800 ;
    RECT 366.660 1.400 367.500 765.800 ;
    RECT 367.780 1.400 368.620 765.800 ;
    RECT 368.900 1.400 369.740 765.800 ;
    RECT 370.020 1.400 370.860 765.800 ;
    RECT 371.140 1.400 371.980 765.800 ;
    RECT 372.260 1.400 373.100 765.800 ;
    RECT 373.380 1.400 374.220 765.800 ;
    RECT 374.500 1.400 375.340 765.800 ;
    RECT 375.620 1.400 376.460 765.800 ;
    RECT 376.740 1.400 377.580 765.800 ;
    RECT 377.860 1.400 378.700 765.800 ;
    RECT 378.980 1.400 379.820 765.800 ;
    RECT 380.100 1.400 380.940 765.800 ;
    RECT 381.220 1.400 382.060 765.800 ;
    RECT 382.340 1.400 383.180 765.800 ;
    RECT 383.460 1.400 384.300 765.800 ;
    RECT 384.580 1.400 385.420 765.800 ;
    RECT 385.700 1.400 386.540 765.800 ;
    RECT 386.820 1.400 387.660 765.800 ;
    RECT 387.940 1.400 388.780 765.800 ;
    RECT 389.060 1.400 389.900 765.800 ;
    RECT 390.180 1.400 391.020 765.800 ;
    RECT 391.300 1.400 392.140 765.800 ;
    RECT 392.420 1.400 393.260 765.800 ;
    RECT 393.540 1.400 394.380 765.800 ;
    RECT 394.660 1.400 395.500 765.800 ;
    RECT 395.780 1.400 396.620 765.800 ;
    RECT 396.900 1.400 397.740 765.800 ;
    RECT 398.020 1.400 398.860 765.800 ;
    RECT 399.140 1.400 399.980 765.800 ;
    RECT 400.260 1.400 401.100 765.800 ;
    RECT 401.380 1.400 402.220 765.800 ;
    RECT 402.500 1.400 403.340 765.800 ;
    RECT 403.620 1.400 404.460 765.800 ;
    RECT 404.740 1.400 405.580 765.800 ;
    RECT 405.860 1.400 406.700 765.800 ;
    RECT 406.980 1.400 407.820 765.800 ;
    RECT 408.100 1.400 408.940 765.800 ;
    RECT 409.220 1.400 410.060 765.800 ;
    RECT 410.340 1.400 411.180 765.800 ;
    RECT 411.460 1.400 412.300 765.800 ;
    RECT 412.580 1.400 413.420 765.800 ;
    RECT 413.700 1.400 414.540 765.800 ;
    RECT 414.820 1.400 415.660 765.800 ;
    RECT 415.940 1.400 416.780 765.800 ;
    RECT 417.060 1.400 417.900 765.800 ;
    RECT 418.180 1.400 419.020 765.800 ;
    RECT 419.300 1.400 420.140 765.800 ;
    RECT 420.420 1.400 421.260 765.800 ;
    RECT 421.540 1.400 422.380 765.800 ;
    RECT 422.660 1.400 423.500 765.800 ;
    RECT 423.780 1.400 424.620 765.800 ;
    RECT 424.900 1.400 425.740 765.800 ;
    RECT 426.020 1.400 426.860 765.800 ;
    RECT 427.140 1.400 427.980 765.800 ;
    RECT 428.260 1.400 429.100 765.800 ;
    RECT 429.380 1.400 430.220 765.800 ;
    RECT 430.500 1.400 431.340 765.800 ;
    RECT 431.620 1.400 432.460 765.800 ;
    RECT 432.740 1.400 433.580 765.800 ;
    RECT 433.860 1.400 434.700 765.800 ;
    RECT 434.980 1.400 435.820 765.800 ;
    RECT 436.100 1.400 436.940 765.800 ;
    RECT 437.220 1.400 438.060 765.800 ;
    RECT 438.340 1.400 439.180 765.800 ;
    RECT 439.460 1.400 440.300 765.800 ;
    RECT 440.580 1.400 441.420 765.800 ;
    RECT 441.700 1.400 442.540 765.800 ;
    RECT 442.820 1.400 443.660 765.800 ;
    RECT 443.940 1.400 444.780 765.800 ;
    RECT 445.060 1.400 445.900 765.800 ;
    RECT 446.180 1.400 447.020 765.800 ;
    RECT 447.300 1.400 448.140 765.800 ;
    RECT 448.420 1.400 449.260 765.800 ;
    RECT 449.540 1.400 450.380 765.800 ;
    RECT 450.660 1.400 451.500 765.800 ;
    RECT 451.780 1.400 452.620 765.800 ;
    RECT 452.900 1.400 453.740 765.800 ;
    RECT 454.020 1.400 454.860 765.800 ;
    RECT 455.140 1.400 455.980 765.800 ;
    RECT 456.260 1.400 457.100 765.800 ;
    RECT 457.380 1.400 458.220 765.800 ;
    RECT 458.500 1.400 459.340 765.800 ;
    RECT 459.620 1.400 460.460 765.800 ;
    RECT 460.740 1.400 461.580 765.800 ;
    RECT 461.860 1.400 462.700 765.800 ;
    RECT 462.980 1.400 463.820 765.800 ;
    RECT 464.100 1.400 464.940 765.800 ;
    RECT 465.220 1.400 466.060 765.800 ;
    RECT 466.340 1.400 467.180 765.800 ;
    RECT 467.460 1.400 468.300 765.800 ;
    RECT 468.580 1.400 469.420 765.800 ;
    RECT 469.700 1.400 470.540 765.800 ;
    RECT 470.820 1.400 471.660 765.800 ;
    RECT 471.940 1.400 472.780 765.800 ;
    RECT 473.060 1.400 473.900 765.800 ;
    RECT 474.180 1.400 475.020 765.800 ;
    RECT 475.300 1.400 476.140 765.800 ;
    RECT 476.420 1.400 477.260 765.800 ;
    RECT 477.540 1.400 478.380 765.800 ;
    RECT 478.660 1.400 479.500 765.800 ;
    RECT 479.780 1.400 480.620 765.800 ;
    RECT 480.900 1.400 481.740 765.800 ;
    RECT 482.020 1.400 482.860 765.800 ;
    RECT 483.140 1.400 483.980 765.800 ;
    RECT 484.260 1.400 485.100 765.800 ;
    RECT 485.380 1.400 486.220 765.800 ;
    RECT 486.500 1.400 487.340 765.800 ;
    RECT 487.620 1.400 488.460 765.800 ;
    RECT 488.740 1.400 489.580 765.800 ;
    RECT 489.860 1.400 490.700 765.800 ;
    RECT 490.980 1.400 491.820 765.800 ;
    RECT 492.100 1.400 492.940 765.800 ;
    RECT 493.220 1.400 494.060 765.800 ;
    RECT 494.340 1.400 495.180 765.800 ;
    RECT 495.460 1.400 496.300 765.800 ;
    RECT 496.580 1.400 497.420 765.800 ;
    RECT 497.700 1.400 498.540 765.800 ;
    RECT 498.820 1.400 499.660 765.800 ;
    RECT 499.940 1.400 500.780 765.800 ;
    RECT 501.060 1.400 501.900 765.800 ;
    RECT 502.180 1.400 503.020 765.800 ;
    RECT 503.300 1.400 504.140 765.800 ;
    RECT 504.420 1.400 505.260 765.800 ;
    RECT 505.540 1.400 506.380 765.800 ;
    RECT 506.660 1.400 507.500 765.800 ;
    RECT 507.780 1.400 508.620 765.800 ;
    RECT 508.900 1.400 509.740 765.800 ;
    RECT 510.020 1.400 510.860 765.800 ;
    RECT 511.140 1.400 511.980 765.800 ;
    RECT 512.260 1.400 513.100 765.800 ;
    RECT 513.380 1.400 514.220 765.800 ;
    RECT 514.500 1.400 515.340 765.800 ;
    RECT 515.620 1.400 516.460 765.800 ;
    RECT 516.740 1.400 517.580 765.800 ;
    RECT 517.860 1.400 518.700 765.800 ;
    RECT 518.980 1.400 519.820 765.800 ;
    RECT 520.100 1.400 520.940 765.800 ;
    RECT 521.220 1.400 522.060 765.800 ;
    RECT 522.340 1.400 523.180 765.800 ;
    RECT 523.460 1.400 524.300 765.800 ;
    RECT 524.580 1.400 525.420 765.800 ;
    RECT 525.700 1.400 526.540 765.800 ;
    RECT 526.820 1.400 527.660 765.800 ;
    RECT 527.940 1.400 528.780 765.800 ;
    RECT 529.060 1.400 529.900 765.800 ;
    RECT 530.180 1.400 531.020 765.800 ;
    RECT 531.300 1.400 532.140 765.800 ;
    RECT 532.420 1.400 533.260 765.800 ;
    RECT 533.540 1.400 534.380 765.800 ;
    RECT 534.660 1.400 535.500 765.800 ;
    RECT 535.780 1.400 536.620 765.800 ;
    RECT 536.900 1.400 537.740 765.800 ;
    RECT 538.020 1.400 538.860 765.800 ;
    RECT 539.140 1.400 539.980 765.800 ;
    RECT 540.260 1.400 541.100 765.800 ;
    RECT 541.380 1.400 542.220 765.800 ;
    RECT 542.500 1.400 543.340 765.800 ;
    RECT 543.620 1.400 544.460 765.800 ;
    RECT 544.740 1.400 545.580 765.800 ;
    RECT 545.860 1.400 546.700 765.800 ;
    RECT 546.980 1.400 547.820 765.800 ;
    RECT 548.100 1.400 548.940 765.800 ;
    RECT 549.220 1.400 550.060 765.800 ;
    RECT 550.340 1.400 551.180 765.800 ;
    RECT 551.460 1.400 552.300 765.800 ;
    RECT 552.580 1.400 553.420 765.800 ;
    RECT 553.700 1.400 554.540 765.800 ;
    RECT 554.820 1.400 555.660 765.800 ;
    RECT 555.940 1.400 556.780 765.800 ;
    RECT 557.060 1.400 557.900 765.800 ;
    RECT 558.180 1.400 559.020 765.800 ;
    RECT 559.300 1.400 560.140 765.800 ;
    RECT 560.420 1.400 561.260 765.800 ;
    RECT 561.540 1.400 562.380 765.800 ;
    RECT 562.660 1.400 563.500 765.800 ;
    RECT 563.780 1.400 564.620 765.800 ;
    RECT 564.900 1.400 565.740 765.800 ;
    RECT 566.020 1.400 566.860 765.800 ;
    RECT 567.140 1.400 567.980 765.800 ;
    RECT 568.260 1.400 569.100 765.800 ;
    RECT 569.380 1.400 570.220 765.800 ;
    RECT 570.500 1.400 571.340 765.800 ;
    RECT 571.620 1.400 572.460 765.800 ;
    RECT 572.740 1.400 573.580 765.800 ;
    RECT 573.860 1.400 574.700 765.800 ;
    RECT 574.980 1.400 575.820 765.800 ;
    RECT 576.100 1.400 576.940 765.800 ;
    RECT 577.220 1.400 578.060 765.800 ;
    RECT 578.340 1.400 579.180 765.800 ;
    RECT 579.460 1.400 580.300 765.800 ;
    RECT 580.580 1.400 581.420 765.800 ;
    RECT 581.700 1.400 582.540 765.800 ;
    RECT 582.820 1.400 583.660 765.800 ;
    RECT 583.940 1.400 584.780 765.800 ;
    RECT 585.060 1.400 585.900 765.800 ;
    RECT 586.180 1.400 587.020 765.800 ;
    RECT 587.300 1.400 588.140 765.800 ;
    RECT 588.420 1.400 589.260 765.800 ;
    RECT 589.540 1.400 590.380 765.800 ;
    RECT 590.660 1.400 591.500 765.800 ;
    RECT 591.780 1.400 592.620 765.800 ;
    RECT 592.900 1.400 593.740 765.800 ;
    RECT 594.020 1.400 594.860 765.800 ;
    RECT 595.140 1.400 595.980 765.800 ;
    RECT 596.260 1.400 597.100 765.800 ;
    RECT 597.380 1.400 598.220 765.800 ;
    RECT 598.500 1.400 599.340 765.800 ;
    RECT 599.620 1.400 600.460 765.800 ;
    RECT 600.740 1.400 601.580 765.800 ;
    RECT 601.860 1.400 602.700 765.800 ;
    RECT 602.980 1.400 603.820 765.800 ;
    RECT 604.100 1.400 604.940 765.800 ;
    RECT 605.220 1.400 606.060 765.800 ;
    RECT 606.340 1.400 607.180 765.800 ;
    RECT 607.460 1.400 608.300 765.800 ;
    RECT 608.580 1.400 609.420 765.800 ;
    RECT 609.700 1.400 610.540 765.800 ;
    RECT 610.820 1.400 611.660 765.800 ;
    RECT 611.940 1.400 612.780 765.800 ;
    RECT 613.060 1.400 613.900 765.800 ;
    RECT 614.180 1.400 615.020 765.800 ;
    RECT 615.300 1.400 616.140 765.800 ;
    RECT 616.420 1.400 617.260 765.800 ;
    RECT 617.540 1.400 618.380 765.800 ;
    RECT 618.660 1.400 619.500 765.800 ;
    RECT 619.780 1.400 620.620 765.800 ;
    RECT 620.900 1.400 621.740 765.800 ;
    RECT 622.020 1.400 622.860 765.800 ;
    RECT 623.140 1.400 623.980 765.800 ;
    RECT 624.260 1.400 625.100 765.800 ;
    RECT 625.380 1.400 626.220 765.800 ;
    RECT 626.500 1.400 627.340 765.800 ;
    RECT 627.620 1.400 628.460 765.800 ;
    RECT 628.740 1.400 629.580 765.800 ;
    RECT 629.860 1.400 630.700 765.800 ;
    RECT 630.980 1.400 631.820 765.800 ;
    RECT 632.100 1.400 632.940 765.800 ;
    RECT 633.220 1.400 634.060 765.800 ;
    RECT 634.340 1.400 635.180 765.800 ;
    RECT 635.460 1.400 636.300 765.800 ;
    RECT 636.580 1.400 637.420 765.800 ;
    RECT 637.700 1.400 638.540 765.800 ;
    RECT 638.820 1.400 639.660 765.800 ;
    RECT 639.940 1.400 640.780 765.800 ;
    RECT 641.060 1.400 641.900 765.800 ;
    RECT 642.180 1.400 643.020 765.800 ;
    RECT 643.300 1.400 644.140 765.800 ;
    RECT 644.420 1.400 645.260 765.800 ;
    RECT 645.540 1.400 646.380 765.800 ;
    RECT 646.660 1.400 647.500 765.800 ;
    RECT 647.780 1.400 648.620 765.800 ;
    RECT 648.900 1.400 649.740 765.800 ;
    RECT 650.020 1.400 650.860 765.800 ;
    RECT 651.140 1.400 651.980 765.800 ;
    RECT 652.260 1.400 653.100 765.800 ;
    RECT 653.380 1.400 654.220 765.800 ;
    RECT 654.500 1.400 655.340 765.800 ;
    RECT 655.620 1.400 656.460 765.800 ;
    RECT 656.740 1.400 657.580 765.800 ;
    RECT 657.860 1.400 658.700 765.800 ;
    RECT 658.980 1.400 659.820 765.800 ;
    RECT 660.100 1.400 660.940 765.800 ;
    RECT 661.220 1.400 662.060 765.800 ;
    RECT 662.340 1.400 663.180 765.800 ;
    RECT 663.460 1.400 664.300 765.800 ;
    RECT 664.580 1.400 665.420 765.800 ;
    RECT 665.700 1.400 666.540 765.800 ;
    RECT 666.820 1.400 667.660 765.800 ;
    RECT 667.940 1.400 668.780 765.800 ;
    RECT 669.060 1.400 669.900 765.800 ;
    RECT 670.180 1.400 671.020 765.800 ;
    RECT 671.300 1.400 672.140 765.800 ;
    RECT 672.420 1.400 673.260 765.800 ;
    RECT 673.540 1.400 674.380 765.800 ;
    RECT 674.660 1.400 675.500 765.800 ;
    RECT 675.780 1.400 676.620 765.800 ;
    RECT 676.900 1.400 677.740 765.800 ;
    RECT 678.020 1.400 678.860 765.800 ;
    RECT 679.140 1.400 679.980 765.800 ;
    RECT 680.260 1.400 681.100 765.800 ;
    RECT 681.380 1.400 682.220 765.800 ;
    RECT 682.500 1.400 683.340 765.800 ;
    RECT 683.620 1.400 684.460 765.800 ;
    RECT 684.740 1.400 685.580 765.800 ;
    RECT 685.860 1.400 686.700 765.800 ;
    RECT 686.980 1.400 689.130 765.800 ;
    LAYER OVERLAP ;
    RECT 0 0 689.130 767.200 ;
  END
END fakeram_512x256_1r1w

END LIBRARY
