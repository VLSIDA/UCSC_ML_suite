VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_1x256_1r1w
  FOREIGN fakeram_1x256_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 130.910 BY 163.800 ;
  CLASS BLOCK ;
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 0.805 0.140 0.875 ;
    END
  END w0_wd_in[0]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1.105 0.000 1.175 0.140 ;
    END
  END r0_rd_out[0]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.725 0.140 18.795 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.645 0.140 36.715 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.140 54.635 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.485 0.140 72.555 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 130.770 0.805 130.910 0.875 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 130.770 18.725 130.910 18.795 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 130.770 36.645 130.910 36.715 ;
    END
  END w0_addr_in[6]
  PIN w0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 130.770 54.565 130.910 54.635 ;
    END
  END w0_addr_in[7]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.405 0.140 90.475 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.325 0.140 108.395 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.245 0.140 126.315 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.165 0.140 144.235 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 130.770 72.485 130.910 72.555 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 130.770 90.405 130.910 90.475 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 130.770 108.325 130.910 108.395 ;
    END
  END r0_addr_in[6]
  PIN r0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 130.770 126.245 130.910 126.315 ;
    END
  END r0_addr_in[7]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1.105 163.660 1.175 163.800 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 22.385 163.660 22.455 163.800 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 43.665 163.660 43.735 163.800 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 64.945 163.660 65.015 163.800 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 86.225 163.660 86.295 163.800 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 0.430 0.700 0.710 163.100 ;
      RECT 2.670 0.700 2.950 163.100 ;
      RECT 4.910 0.700 5.190 163.100 ;
      RECT 7.150 0.700 7.430 163.100 ;
      RECT 9.390 0.700 9.670 163.100 ;
      RECT 11.630 0.700 11.910 163.100 ;
      RECT 13.870 0.700 14.150 163.100 ;
      RECT 16.110 0.700 16.390 163.100 ;
      RECT 18.350 0.700 18.630 163.100 ;
      RECT 20.590 0.700 20.870 163.100 ;
      RECT 22.830 0.700 23.110 163.100 ;
      RECT 25.070 0.700 25.350 163.100 ;
      RECT 27.310 0.700 27.590 163.100 ;
      RECT 29.550 0.700 29.830 163.100 ;
      RECT 31.790 0.700 32.070 163.100 ;
      RECT 34.030 0.700 34.310 163.100 ;
      RECT 36.270 0.700 36.550 163.100 ;
      RECT 38.510 0.700 38.790 163.100 ;
      RECT 40.750 0.700 41.030 163.100 ;
      RECT 42.990 0.700 43.270 163.100 ;
      RECT 45.230 0.700 45.510 163.100 ;
      RECT 47.470 0.700 47.750 163.100 ;
      RECT 49.710 0.700 49.990 163.100 ;
      RECT 51.950 0.700 52.230 163.100 ;
      RECT 54.190 0.700 54.470 163.100 ;
      RECT 56.430 0.700 56.710 163.100 ;
      RECT 58.670 0.700 58.950 163.100 ;
      RECT 60.910 0.700 61.190 163.100 ;
      RECT 63.150 0.700 63.430 163.100 ;
      RECT 65.390 0.700 65.670 163.100 ;
      RECT 67.630 0.700 67.910 163.100 ;
      RECT 69.870 0.700 70.150 163.100 ;
      RECT 72.110 0.700 72.390 163.100 ;
      RECT 74.350 0.700 74.630 163.100 ;
      RECT 76.590 0.700 76.870 163.100 ;
      RECT 78.830 0.700 79.110 163.100 ;
      RECT 81.070 0.700 81.350 163.100 ;
      RECT 83.310 0.700 83.590 163.100 ;
      RECT 85.550 0.700 85.830 163.100 ;
      RECT 87.790 0.700 88.070 163.100 ;
      RECT 90.030 0.700 90.310 163.100 ;
      RECT 92.270 0.700 92.550 163.100 ;
      RECT 94.510 0.700 94.790 163.100 ;
      RECT 96.750 0.700 97.030 163.100 ;
      RECT 98.990 0.700 99.270 163.100 ;
      RECT 101.230 0.700 101.510 163.100 ;
      RECT 103.470 0.700 103.750 163.100 ;
      RECT 105.710 0.700 105.990 163.100 ;
      RECT 107.950 0.700 108.230 163.100 ;
      RECT 110.190 0.700 110.470 163.100 ;
      RECT 112.430 0.700 112.710 163.100 ;
      RECT 114.670 0.700 114.950 163.100 ;
      RECT 116.910 0.700 117.190 163.100 ;
      RECT 119.150 0.700 119.430 163.100 ;
      RECT 121.390 0.700 121.670 163.100 ;
      RECT 123.630 0.700 123.910 163.100 ;
      RECT 125.870 0.700 126.150 163.100 ;
      RECT 128.110 0.700 128.390 163.100 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 0.430 0.700 0.710 163.100 ;
      RECT 2.670 0.700 2.950 163.100 ;
      RECT 4.910 0.700 5.190 163.100 ;
      RECT 7.150 0.700 7.430 163.100 ;
      RECT 9.390 0.700 9.670 163.100 ;
      RECT 11.630 0.700 11.910 163.100 ;
      RECT 13.870 0.700 14.150 163.100 ;
      RECT 16.110 0.700 16.390 163.100 ;
      RECT 18.350 0.700 18.630 163.100 ;
      RECT 20.590 0.700 20.870 163.100 ;
      RECT 22.830 0.700 23.110 163.100 ;
      RECT 25.070 0.700 25.350 163.100 ;
      RECT 27.310 0.700 27.590 163.100 ;
      RECT 29.550 0.700 29.830 163.100 ;
      RECT 31.790 0.700 32.070 163.100 ;
      RECT 34.030 0.700 34.310 163.100 ;
      RECT 36.270 0.700 36.550 163.100 ;
      RECT 38.510 0.700 38.790 163.100 ;
      RECT 40.750 0.700 41.030 163.100 ;
      RECT 42.990 0.700 43.270 163.100 ;
      RECT 45.230 0.700 45.510 163.100 ;
      RECT 47.470 0.700 47.750 163.100 ;
      RECT 49.710 0.700 49.990 163.100 ;
      RECT 51.950 0.700 52.230 163.100 ;
      RECT 54.190 0.700 54.470 163.100 ;
      RECT 56.430 0.700 56.710 163.100 ;
      RECT 58.670 0.700 58.950 163.100 ;
      RECT 60.910 0.700 61.190 163.100 ;
      RECT 63.150 0.700 63.430 163.100 ;
      RECT 65.390 0.700 65.670 163.100 ;
      RECT 67.630 0.700 67.910 163.100 ;
      RECT 69.870 0.700 70.150 163.100 ;
      RECT 72.110 0.700 72.390 163.100 ;
      RECT 74.350 0.700 74.630 163.100 ;
      RECT 76.590 0.700 76.870 163.100 ;
      RECT 78.830 0.700 79.110 163.100 ;
      RECT 81.070 0.700 81.350 163.100 ;
      RECT 83.310 0.700 83.590 163.100 ;
      RECT 85.550 0.700 85.830 163.100 ;
      RECT 87.790 0.700 88.070 163.100 ;
      RECT 90.030 0.700 90.310 163.100 ;
      RECT 92.270 0.700 92.550 163.100 ;
      RECT 94.510 0.700 94.790 163.100 ;
      RECT 96.750 0.700 97.030 163.100 ;
      RECT 98.990 0.700 99.270 163.100 ;
      RECT 101.230 0.700 101.510 163.100 ;
      RECT 103.470 0.700 103.750 163.100 ;
      RECT 105.710 0.700 105.990 163.100 ;
      RECT 107.950 0.700 108.230 163.100 ;
      RECT 110.190 0.700 110.470 163.100 ;
      RECT 112.430 0.700 112.710 163.100 ;
      RECT 114.670 0.700 114.950 163.100 ;
      RECT 116.910 0.700 117.190 163.100 ;
      RECT 119.150 0.700 119.430 163.100 ;
      RECT 121.390 0.700 121.670 163.100 ;
      RECT 123.630 0.700 123.910 163.100 ;
      RECT 125.870 0.700 126.150 163.100 ;
      RECT 128.110 0.700 128.390 163.100 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 130.910 163.800 ;
    LAYER metal2 ;
    RECT 0 0 130.910 163.800 ;
    LAYER metal3 ;
    RECT 0 0 130.910 163.800 ;
    LAYER metal4 ;
    RECT 0 0 130.910 163.800 ;
    LAYER OVERLAP ;
    RECT 0 0 130.910 163.800 ;
  END
END fakeram_1x256_1r1w

END LIBRARY
