VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_512x2048_1r1w
  FOREIGN fakeram_512x2048_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 5871.900 BY 1436.160 ;
  CLASS BLOCK ;
  PIN w0_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 6.650 0.800 6.950 ;
    END
  END w0_mask_in[0]
  PIN w0_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 8.010 0.800 8.310 ;
    END
  END w0_mask_in[1]
  PIN w0_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 9.370 0.800 9.670 ;
    END
  END w0_mask_in[2]
  PIN w0_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 10.730 0.800 11.030 ;
    END
  END w0_mask_in[3]
  PIN w0_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 12.090 0.800 12.390 ;
    END
  END w0_mask_in[4]
  PIN w0_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 13.450 0.800 13.750 ;
    END
  END w0_mask_in[5]
  PIN w0_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.810 0.800 15.110 ;
    END
  END w0_mask_in[6]
  PIN w0_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 16.170 0.800 16.470 ;
    END
  END w0_mask_in[7]
  PIN w0_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 17.530 0.800 17.830 ;
    END
  END w0_mask_in[8]
  PIN w0_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 18.890 0.800 19.190 ;
    END
  END w0_mask_in[9]
  PIN w0_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.250 0.800 20.550 ;
    END
  END w0_mask_in[10]
  PIN w0_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 21.610 0.800 21.910 ;
    END
  END w0_mask_in[11]
  PIN w0_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.970 0.800 23.270 ;
    END
  END w0_mask_in[12]
  PIN w0_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 24.330 0.800 24.630 ;
    END
  END w0_mask_in[13]
  PIN w0_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 25.690 0.800 25.990 ;
    END
  END w0_mask_in[14]
  PIN w0_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 27.050 0.800 27.350 ;
    END
  END w0_mask_in[15]
  PIN w0_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 28.410 0.800 28.710 ;
    END
  END w0_mask_in[16]
  PIN w0_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 29.770 0.800 30.070 ;
    END
  END w0_mask_in[17]
  PIN w0_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.130 0.800 31.430 ;
    END
  END w0_mask_in[18]
  PIN w0_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 32.490 0.800 32.790 ;
    END
  END w0_mask_in[19]
  PIN w0_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 33.850 0.800 34.150 ;
    END
  END w0_mask_in[20]
  PIN w0_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 35.210 0.800 35.510 ;
    END
  END w0_mask_in[21]
  PIN w0_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 36.570 0.800 36.870 ;
    END
  END w0_mask_in[22]
  PIN w0_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.930 0.800 38.230 ;
    END
  END w0_mask_in[23]
  PIN w0_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.290 0.800 39.590 ;
    END
  END w0_mask_in[24]
  PIN w0_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.650 0.800 40.950 ;
    END
  END w0_mask_in[25]
  PIN w0_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 42.010 0.800 42.310 ;
    END
  END w0_mask_in[26]
  PIN w0_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 43.370 0.800 43.670 ;
    END
  END w0_mask_in[27]
  PIN w0_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 44.730 0.800 45.030 ;
    END
  END w0_mask_in[28]
  PIN w0_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 46.090 0.800 46.390 ;
    END
  END w0_mask_in[29]
  PIN w0_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 47.450 0.800 47.750 ;
    END
  END w0_mask_in[30]
  PIN w0_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 48.810 0.800 49.110 ;
    END
  END w0_mask_in[31]
  PIN w0_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 50.170 0.800 50.470 ;
    END
  END w0_mask_in[32]
  PIN w0_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 51.530 0.800 51.830 ;
    END
  END w0_mask_in[33]
  PIN w0_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 52.890 0.800 53.190 ;
    END
  END w0_mask_in[34]
  PIN w0_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 54.250 0.800 54.550 ;
    END
  END w0_mask_in[35]
  PIN w0_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.610 0.800 55.910 ;
    END
  END w0_mask_in[36]
  PIN w0_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 56.970 0.800 57.270 ;
    END
  END w0_mask_in[37]
  PIN w0_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 58.330 0.800 58.630 ;
    END
  END w0_mask_in[38]
  PIN w0_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 59.690 0.800 59.990 ;
    END
  END w0_mask_in[39]
  PIN w0_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 61.050 0.800 61.350 ;
    END
  END w0_mask_in[40]
  PIN w0_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 62.410 0.800 62.710 ;
    END
  END w0_mask_in[41]
  PIN w0_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 63.770 0.800 64.070 ;
    END
  END w0_mask_in[42]
  PIN w0_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 65.130 0.800 65.430 ;
    END
  END w0_mask_in[43]
  PIN w0_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 66.490 0.800 66.790 ;
    END
  END w0_mask_in[44]
  PIN w0_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.850 0.800 68.150 ;
    END
  END w0_mask_in[45]
  PIN w0_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 69.210 0.800 69.510 ;
    END
  END w0_mask_in[46]
  PIN w0_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 70.570 0.800 70.870 ;
    END
  END w0_mask_in[47]
  PIN w0_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.930 0.800 72.230 ;
    END
  END w0_mask_in[48]
  PIN w0_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 73.290 0.800 73.590 ;
    END
  END w0_mask_in[49]
  PIN w0_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 74.650 0.800 74.950 ;
    END
  END w0_mask_in[50]
  PIN w0_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.010 0.800 76.310 ;
    END
  END w0_mask_in[51]
  PIN w0_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 77.370 0.800 77.670 ;
    END
  END w0_mask_in[52]
  PIN w0_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 78.730 0.800 79.030 ;
    END
  END w0_mask_in[53]
  PIN w0_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 80.090 0.800 80.390 ;
    END
  END w0_mask_in[54]
  PIN w0_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 81.450 0.800 81.750 ;
    END
  END w0_mask_in[55]
  PIN w0_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 82.810 0.800 83.110 ;
    END
  END w0_mask_in[56]
  PIN w0_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 84.170 0.800 84.470 ;
    END
  END w0_mask_in[57]
  PIN w0_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 85.530 0.800 85.830 ;
    END
  END w0_mask_in[58]
  PIN w0_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 86.890 0.800 87.190 ;
    END
  END w0_mask_in[59]
  PIN w0_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 88.250 0.800 88.550 ;
    END
  END w0_mask_in[60]
  PIN w0_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.610 0.800 89.910 ;
    END
  END w0_mask_in[61]
  PIN w0_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 90.970 0.800 91.270 ;
    END
  END w0_mask_in[62]
  PIN w0_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 92.330 0.800 92.630 ;
    END
  END w0_mask_in[63]
  PIN w0_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 93.690 0.800 93.990 ;
    END
  END w0_mask_in[64]
  PIN w0_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 95.050 0.800 95.350 ;
    END
  END w0_mask_in[65]
  PIN w0_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 96.410 0.800 96.710 ;
    END
  END w0_mask_in[66]
  PIN w0_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 97.770 0.800 98.070 ;
    END
  END w0_mask_in[67]
  PIN w0_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 99.130 0.800 99.430 ;
    END
  END w0_mask_in[68]
  PIN w0_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 100.490 0.800 100.790 ;
    END
  END w0_mask_in[69]
  PIN w0_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 101.850 0.800 102.150 ;
    END
  END w0_mask_in[70]
  PIN w0_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 103.210 0.800 103.510 ;
    END
  END w0_mask_in[71]
  PIN w0_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 104.570 0.800 104.870 ;
    END
  END w0_mask_in[72]
  PIN w0_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 105.930 0.800 106.230 ;
    END
  END w0_mask_in[73]
  PIN w0_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 107.290 0.800 107.590 ;
    END
  END w0_mask_in[74]
  PIN w0_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 108.650 0.800 108.950 ;
    END
  END w0_mask_in[75]
  PIN w0_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 110.010 0.800 110.310 ;
    END
  END w0_mask_in[76]
  PIN w0_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 111.370 0.800 111.670 ;
    END
  END w0_mask_in[77]
  PIN w0_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 112.730 0.800 113.030 ;
    END
  END w0_mask_in[78]
  PIN w0_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 114.090 0.800 114.390 ;
    END
  END w0_mask_in[79]
  PIN w0_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 115.450 0.800 115.750 ;
    END
  END w0_mask_in[80]
  PIN w0_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 116.810 0.800 117.110 ;
    END
  END w0_mask_in[81]
  PIN w0_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 118.170 0.800 118.470 ;
    END
  END w0_mask_in[82]
  PIN w0_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 119.530 0.800 119.830 ;
    END
  END w0_mask_in[83]
  PIN w0_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 120.890 0.800 121.190 ;
    END
  END w0_mask_in[84]
  PIN w0_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 122.250 0.800 122.550 ;
    END
  END w0_mask_in[85]
  PIN w0_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 123.610 0.800 123.910 ;
    END
  END w0_mask_in[86]
  PIN w0_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 124.970 0.800 125.270 ;
    END
  END w0_mask_in[87]
  PIN w0_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 126.330 0.800 126.630 ;
    END
  END w0_mask_in[88]
  PIN w0_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 127.690 0.800 127.990 ;
    END
  END w0_mask_in[89]
  PIN w0_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 129.050 0.800 129.350 ;
    END
  END w0_mask_in[90]
  PIN w0_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 130.410 0.800 130.710 ;
    END
  END w0_mask_in[91]
  PIN w0_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 131.770 0.800 132.070 ;
    END
  END w0_mask_in[92]
  PIN w0_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 133.130 0.800 133.430 ;
    END
  END w0_mask_in[93]
  PIN w0_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 134.490 0.800 134.790 ;
    END
  END w0_mask_in[94]
  PIN w0_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 135.850 0.800 136.150 ;
    END
  END w0_mask_in[95]
  PIN w0_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 137.210 0.800 137.510 ;
    END
  END w0_mask_in[96]
  PIN w0_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 138.570 0.800 138.870 ;
    END
  END w0_mask_in[97]
  PIN w0_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.930 0.800 140.230 ;
    END
  END w0_mask_in[98]
  PIN w0_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 141.290 0.800 141.590 ;
    END
  END w0_mask_in[99]
  PIN w0_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 142.650 0.800 142.950 ;
    END
  END w0_mask_in[100]
  PIN w0_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 144.010 0.800 144.310 ;
    END
  END w0_mask_in[101]
  PIN w0_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 145.370 0.800 145.670 ;
    END
  END w0_mask_in[102]
  PIN w0_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 146.730 0.800 147.030 ;
    END
  END w0_mask_in[103]
  PIN w0_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 148.090 0.800 148.390 ;
    END
  END w0_mask_in[104]
  PIN w0_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 149.450 0.800 149.750 ;
    END
  END w0_mask_in[105]
  PIN w0_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 150.810 0.800 151.110 ;
    END
  END w0_mask_in[106]
  PIN w0_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 152.170 0.800 152.470 ;
    END
  END w0_mask_in[107]
  PIN w0_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 153.530 0.800 153.830 ;
    END
  END w0_mask_in[108]
  PIN w0_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 154.890 0.800 155.190 ;
    END
  END w0_mask_in[109]
  PIN w0_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 156.250 0.800 156.550 ;
    END
  END w0_mask_in[110]
  PIN w0_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 157.610 0.800 157.910 ;
    END
  END w0_mask_in[111]
  PIN w0_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 158.970 0.800 159.270 ;
    END
  END w0_mask_in[112]
  PIN w0_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 160.330 0.800 160.630 ;
    END
  END w0_mask_in[113]
  PIN w0_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 161.690 0.800 161.990 ;
    END
  END w0_mask_in[114]
  PIN w0_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 163.050 0.800 163.350 ;
    END
  END w0_mask_in[115]
  PIN w0_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 164.410 0.800 164.710 ;
    END
  END w0_mask_in[116]
  PIN w0_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 165.770 0.800 166.070 ;
    END
  END w0_mask_in[117]
  PIN w0_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 167.130 0.800 167.430 ;
    END
  END w0_mask_in[118]
  PIN w0_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 168.490 0.800 168.790 ;
    END
  END w0_mask_in[119]
  PIN w0_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 169.850 0.800 170.150 ;
    END
  END w0_mask_in[120]
  PIN w0_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 171.210 0.800 171.510 ;
    END
  END w0_mask_in[121]
  PIN w0_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 172.570 0.800 172.870 ;
    END
  END w0_mask_in[122]
  PIN w0_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 173.930 0.800 174.230 ;
    END
  END w0_mask_in[123]
  PIN w0_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 175.290 0.800 175.590 ;
    END
  END w0_mask_in[124]
  PIN w0_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 176.650 0.800 176.950 ;
    END
  END w0_mask_in[125]
  PIN w0_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 178.010 0.800 178.310 ;
    END
  END w0_mask_in[126]
  PIN w0_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 179.370 0.800 179.670 ;
    END
  END w0_mask_in[127]
  PIN w0_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 180.730 0.800 181.030 ;
    END
  END w0_mask_in[128]
  PIN w0_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 182.090 0.800 182.390 ;
    END
  END w0_mask_in[129]
  PIN w0_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 183.450 0.800 183.750 ;
    END
  END w0_mask_in[130]
  PIN w0_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 184.810 0.800 185.110 ;
    END
  END w0_mask_in[131]
  PIN w0_mask_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 186.170 0.800 186.470 ;
    END
  END w0_mask_in[132]
  PIN w0_mask_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 187.530 0.800 187.830 ;
    END
  END w0_mask_in[133]
  PIN w0_mask_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 188.890 0.800 189.190 ;
    END
  END w0_mask_in[134]
  PIN w0_mask_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 190.250 0.800 190.550 ;
    END
  END w0_mask_in[135]
  PIN w0_mask_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 191.610 0.800 191.910 ;
    END
  END w0_mask_in[136]
  PIN w0_mask_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 192.970 0.800 193.270 ;
    END
  END w0_mask_in[137]
  PIN w0_mask_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 194.330 0.800 194.630 ;
    END
  END w0_mask_in[138]
  PIN w0_mask_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 195.690 0.800 195.990 ;
    END
  END w0_mask_in[139]
  PIN w0_mask_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 197.050 0.800 197.350 ;
    END
  END w0_mask_in[140]
  PIN w0_mask_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 198.410 0.800 198.710 ;
    END
  END w0_mask_in[141]
  PIN w0_mask_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 199.770 0.800 200.070 ;
    END
  END w0_mask_in[142]
  PIN w0_mask_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 201.130 0.800 201.430 ;
    END
  END w0_mask_in[143]
  PIN w0_mask_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 202.490 0.800 202.790 ;
    END
  END w0_mask_in[144]
  PIN w0_mask_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 203.850 0.800 204.150 ;
    END
  END w0_mask_in[145]
  PIN w0_mask_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 205.210 0.800 205.510 ;
    END
  END w0_mask_in[146]
  PIN w0_mask_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 206.570 0.800 206.870 ;
    END
  END w0_mask_in[147]
  PIN w0_mask_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 207.930 0.800 208.230 ;
    END
  END w0_mask_in[148]
  PIN w0_mask_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 209.290 0.800 209.590 ;
    END
  END w0_mask_in[149]
  PIN w0_mask_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 210.650 0.800 210.950 ;
    END
  END w0_mask_in[150]
  PIN w0_mask_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 212.010 0.800 212.310 ;
    END
  END w0_mask_in[151]
  PIN w0_mask_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 213.370 0.800 213.670 ;
    END
  END w0_mask_in[152]
  PIN w0_mask_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 214.730 0.800 215.030 ;
    END
  END w0_mask_in[153]
  PIN w0_mask_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 216.090 0.800 216.390 ;
    END
  END w0_mask_in[154]
  PIN w0_mask_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 217.450 0.800 217.750 ;
    END
  END w0_mask_in[155]
  PIN w0_mask_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 218.810 0.800 219.110 ;
    END
  END w0_mask_in[156]
  PIN w0_mask_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 220.170 0.800 220.470 ;
    END
  END w0_mask_in[157]
  PIN w0_mask_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 221.530 0.800 221.830 ;
    END
  END w0_mask_in[158]
  PIN w0_mask_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 222.890 0.800 223.190 ;
    END
  END w0_mask_in[159]
  PIN w0_mask_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 224.250 0.800 224.550 ;
    END
  END w0_mask_in[160]
  PIN w0_mask_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 225.610 0.800 225.910 ;
    END
  END w0_mask_in[161]
  PIN w0_mask_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 226.970 0.800 227.270 ;
    END
  END w0_mask_in[162]
  PIN w0_mask_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 228.330 0.800 228.630 ;
    END
  END w0_mask_in[163]
  PIN w0_mask_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 229.690 0.800 229.990 ;
    END
  END w0_mask_in[164]
  PIN w0_mask_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 231.050 0.800 231.350 ;
    END
  END w0_mask_in[165]
  PIN w0_mask_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 232.410 0.800 232.710 ;
    END
  END w0_mask_in[166]
  PIN w0_mask_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 233.770 0.800 234.070 ;
    END
  END w0_mask_in[167]
  PIN w0_mask_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 235.130 0.800 235.430 ;
    END
  END w0_mask_in[168]
  PIN w0_mask_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 236.490 0.800 236.790 ;
    END
  END w0_mask_in[169]
  PIN w0_mask_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 237.850 0.800 238.150 ;
    END
  END w0_mask_in[170]
  PIN w0_mask_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 239.210 0.800 239.510 ;
    END
  END w0_mask_in[171]
  PIN w0_mask_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 240.570 0.800 240.870 ;
    END
  END w0_mask_in[172]
  PIN w0_mask_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 241.930 0.800 242.230 ;
    END
  END w0_mask_in[173]
  PIN w0_mask_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 243.290 0.800 243.590 ;
    END
  END w0_mask_in[174]
  PIN w0_mask_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 244.650 0.800 244.950 ;
    END
  END w0_mask_in[175]
  PIN w0_mask_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 246.010 0.800 246.310 ;
    END
  END w0_mask_in[176]
  PIN w0_mask_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 247.370 0.800 247.670 ;
    END
  END w0_mask_in[177]
  PIN w0_mask_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 248.730 0.800 249.030 ;
    END
  END w0_mask_in[178]
  PIN w0_mask_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 250.090 0.800 250.390 ;
    END
  END w0_mask_in[179]
  PIN w0_mask_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 251.450 0.800 251.750 ;
    END
  END w0_mask_in[180]
  PIN w0_mask_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 252.810 0.800 253.110 ;
    END
  END w0_mask_in[181]
  PIN w0_mask_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 254.170 0.800 254.470 ;
    END
  END w0_mask_in[182]
  PIN w0_mask_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 255.530 0.800 255.830 ;
    END
  END w0_mask_in[183]
  PIN w0_mask_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 256.890 0.800 257.190 ;
    END
  END w0_mask_in[184]
  PIN w0_mask_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 258.250 0.800 258.550 ;
    END
  END w0_mask_in[185]
  PIN w0_mask_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 259.610 0.800 259.910 ;
    END
  END w0_mask_in[186]
  PIN w0_mask_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 260.970 0.800 261.270 ;
    END
  END w0_mask_in[187]
  PIN w0_mask_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 262.330 0.800 262.630 ;
    END
  END w0_mask_in[188]
  PIN w0_mask_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 263.690 0.800 263.990 ;
    END
  END w0_mask_in[189]
  PIN w0_mask_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 265.050 0.800 265.350 ;
    END
  END w0_mask_in[190]
  PIN w0_mask_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 266.410 0.800 266.710 ;
    END
  END w0_mask_in[191]
  PIN w0_mask_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 267.770 0.800 268.070 ;
    END
  END w0_mask_in[192]
  PIN w0_mask_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 269.130 0.800 269.430 ;
    END
  END w0_mask_in[193]
  PIN w0_mask_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 270.490 0.800 270.790 ;
    END
  END w0_mask_in[194]
  PIN w0_mask_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 271.850 0.800 272.150 ;
    END
  END w0_mask_in[195]
  PIN w0_mask_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 273.210 0.800 273.510 ;
    END
  END w0_mask_in[196]
  PIN w0_mask_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 274.570 0.800 274.870 ;
    END
  END w0_mask_in[197]
  PIN w0_mask_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 275.930 0.800 276.230 ;
    END
  END w0_mask_in[198]
  PIN w0_mask_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 277.290 0.800 277.590 ;
    END
  END w0_mask_in[199]
  PIN w0_mask_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 278.650 0.800 278.950 ;
    END
  END w0_mask_in[200]
  PIN w0_mask_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 280.010 0.800 280.310 ;
    END
  END w0_mask_in[201]
  PIN w0_mask_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 281.370 0.800 281.670 ;
    END
  END w0_mask_in[202]
  PIN w0_mask_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 282.730 0.800 283.030 ;
    END
  END w0_mask_in[203]
  PIN w0_mask_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 284.090 0.800 284.390 ;
    END
  END w0_mask_in[204]
  PIN w0_mask_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 285.450 0.800 285.750 ;
    END
  END w0_mask_in[205]
  PIN w0_mask_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 286.810 0.800 287.110 ;
    END
  END w0_mask_in[206]
  PIN w0_mask_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 288.170 0.800 288.470 ;
    END
  END w0_mask_in[207]
  PIN w0_mask_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 289.530 0.800 289.830 ;
    END
  END w0_mask_in[208]
  PIN w0_mask_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 290.890 0.800 291.190 ;
    END
  END w0_mask_in[209]
  PIN w0_mask_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 292.250 0.800 292.550 ;
    END
  END w0_mask_in[210]
  PIN w0_mask_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 293.610 0.800 293.910 ;
    END
  END w0_mask_in[211]
  PIN w0_mask_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 294.970 0.800 295.270 ;
    END
  END w0_mask_in[212]
  PIN w0_mask_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 296.330 0.800 296.630 ;
    END
  END w0_mask_in[213]
  PIN w0_mask_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 297.690 0.800 297.990 ;
    END
  END w0_mask_in[214]
  PIN w0_mask_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 299.050 0.800 299.350 ;
    END
  END w0_mask_in[215]
  PIN w0_mask_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 300.410 0.800 300.710 ;
    END
  END w0_mask_in[216]
  PIN w0_mask_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 301.770 0.800 302.070 ;
    END
  END w0_mask_in[217]
  PIN w0_mask_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 303.130 0.800 303.430 ;
    END
  END w0_mask_in[218]
  PIN w0_mask_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 304.490 0.800 304.790 ;
    END
  END w0_mask_in[219]
  PIN w0_mask_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 305.850 0.800 306.150 ;
    END
  END w0_mask_in[220]
  PIN w0_mask_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 307.210 0.800 307.510 ;
    END
  END w0_mask_in[221]
  PIN w0_mask_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 308.570 0.800 308.870 ;
    END
  END w0_mask_in[222]
  PIN w0_mask_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 309.930 0.800 310.230 ;
    END
  END w0_mask_in[223]
  PIN w0_mask_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 311.290 0.800 311.590 ;
    END
  END w0_mask_in[224]
  PIN w0_mask_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 312.650 0.800 312.950 ;
    END
  END w0_mask_in[225]
  PIN w0_mask_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 314.010 0.800 314.310 ;
    END
  END w0_mask_in[226]
  PIN w0_mask_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 315.370 0.800 315.670 ;
    END
  END w0_mask_in[227]
  PIN w0_mask_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 316.730 0.800 317.030 ;
    END
  END w0_mask_in[228]
  PIN w0_mask_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 318.090 0.800 318.390 ;
    END
  END w0_mask_in[229]
  PIN w0_mask_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 319.450 0.800 319.750 ;
    END
  END w0_mask_in[230]
  PIN w0_mask_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 320.810 0.800 321.110 ;
    END
  END w0_mask_in[231]
  PIN w0_mask_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 322.170 0.800 322.470 ;
    END
  END w0_mask_in[232]
  PIN w0_mask_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 323.530 0.800 323.830 ;
    END
  END w0_mask_in[233]
  PIN w0_mask_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 324.890 0.800 325.190 ;
    END
  END w0_mask_in[234]
  PIN w0_mask_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 326.250 0.800 326.550 ;
    END
  END w0_mask_in[235]
  PIN w0_mask_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 327.610 0.800 327.910 ;
    END
  END w0_mask_in[236]
  PIN w0_mask_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 328.970 0.800 329.270 ;
    END
  END w0_mask_in[237]
  PIN w0_mask_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 330.330 0.800 330.630 ;
    END
  END w0_mask_in[238]
  PIN w0_mask_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 331.690 0.800 331.990 ;
    END
  END w0_mask_in[239]
  PIN w0_mask_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 333.050 0.800 333.350 ;
    END
  END w0_mask_in[240]
  PIN w0_mask_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 334.410 0.800 334.710 ;
    END
  END w0_mask_in[241]
  PIN w0_mask_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 335.770 0.800 336.070 ;
    END
  END w0_mask_in[242]
  PIN w0_mask_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 337.130 0.800 337.430 ;
    END
  END w0_mask_in[243]
  PIN w0_mask_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 338.490 0.800 338.790 ;
    END
  END w0_mask_in[244]
  PIN w0_mask_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 339.850 0.800 340.150 ;
    END
  END w0_mask_in[245]
  PIN w0_mask_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 341.210 0.800 341.510 ;
    END
  END w0_mask_in[246]
  PIN w0_mask_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 342.570 0.800 342.870 ;
    END
  END w0_mask_in[247]
  PIN w0_mask_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 343.930 0.800 344.230 ;
    END
  END w0_mask_in[248]
  PIN w0_mask_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 345.290 0.800 345.590 ;
    END
  END w0_mask_in[249]
  PIN w0_mask_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 346.650 0.800 346.950 ;
    END
  END w0_mask_in[250]
  PIN w0_mask_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 348.010 0.800 348.310 ;
    END
  END w0_mask_in[251]
  PIN w0_mask_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 349.370 0.800 349.670 ;
    END
  END w0_mask_in[252]
  PIN w0_mask_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 350.730 0.800 351.030 ;
    END
  END w0_mask_in[253]
  PIN w0_mask_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 352.090 0.800 352.390 ;
    END
  END w0_mask_in[254]
  PIN w0_mask_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 353.450 0.800 353.750 ;
    END
  END w0_mask_in[255]
  PIN w0_mask_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 354.810 0.800 355.110 ;
    END
  END w0_mask_in[256]
  PIN w0_mask_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 356.170 0.800 356.470 ;
    END
  END w0_mask_in[257]
  PIN w0_mask_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 357.530 0.800 357.830 ;
    END
  END w0_mask_in[258]
  PIN w0_mask_in[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 358.890 0.800 359.190 ;
    END
  END w0_mask_in[259]
  PIN w0_mask_in[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 360.250 0.800 360.550 ;
    END
  END w0_mask_in[260]
  PIN w0_mask_in[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 361.610 0.800 361.910 ;
    END
  END w0_mask_in[261]
  PIN w0_mask_in[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 362.970 0.800 363.270 ;
    END
  END w0_mask_in[262]
  PIN w0_mask_in[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 364.330 0.800 364.630 ;
    END
  END w0_mask_in[263]
  PIN w0_mask_in[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 365.690 0.800 365.990 ;
    END
  END w0_mask_in[264]
  PIN w0_mask_in[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 367.050 0.800 367.350 ;
    END
  END w0_mask_in[265]
  PIN w0_mask_in[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 368.410 0.800 368.710 ;
    END
  END w0_mask_in[266]
  PIN w0_mask_in[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 369.770 0.800 370.070 ;
    END
  END w0_mask_in[267]
  PIN w0_mask_in[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 371.130 0.800 371.430 ;
    END
  END w0_mask_in[268]
  PIN w0_mask_in[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 372.490 0.800 372.790 ;
    END
  END w0_mask_in[269]
  PIN w0_mask_in[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 373.850 0.800 374.150 ;
    END
  END w0_mask_in[270]
  PIN w0_mask_in[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 375.210 0.800 375.510 ;
    END
  END w0_mask_in[271]
  PIN w0_mask_in[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 376.570 0.800 376.870 ;
    END
  END w0_mask_in[272]
  PIN w0_mask_in[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 377.930 0.800 378.230 ;
    END
  END w0_mask_in[273]
  PIN w0_mask_in[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 379.290 0.800 379.590 ;
    END
  END w0_mask_in[274]
  PIN w0_mask_in[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 380.650 0.800 380.950 ;
    END
  END w0_mask_in[275]
  PIN w0_mask_in[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 382.010 0.800 382.310 ;
    END
  END w0_mask_in[276]
  PIN w0_mask_in[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 383.370 0.800 383.670 ;
    END
  END w0_mask_in[277]
  PIN w0_mask_in[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 384.730 0.800 385.030 ;
    END
  END w0_mask_in[278]
  PIN w0_mask_in[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 386.090 0.800 386.390 ;
    END
  END w0_mask_in[279]
  PIN w0_mask_in[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 387.450 0.800 387.750 ;
    END
  END w0_mask_in[280]
  PIN w0_mask_in[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 388.810 0.800 389.110 ;
    END
  END w0_mask_in[281]
  PIN w0_mask_in[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 390.170 0.800 390.470 ;
    END
  END w0_mask_in[282]
  PIN w0_mask_in[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 391.530 0.800 391.830 ;
    END
  END w0_mask_in[283]
  PIN w0_mask_in[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 392.890 0.800 393.190 ;
    END
  END w0_mask_in[284]
  PIN w0_mask_in[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 394.250 0.800 394.550 ;
    END
  END w0_mask_in[285]
  PIN w0_mask_in[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 395.610 0.800 395.910 ;
    END
  END w0_mask_in[286]
  PIN w0_mask_in[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 396.970 0.800 397.270 ;
    END
  END w0_mask_in[287]
  PIN w0_mask_in[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 398.330 0.800 398.630 ;
    END
  END w0_mask_in[288]
  PIN w0_mask_in[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 399.690 0.800 399.990 ;
    END
  END w0_mask_in[289]
  PIN w0_mask_in[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 401.050 0.800 401.350 ;
    END
  END w0_mask_in[290]
  PIN w0_mask_in[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 402.410 0.800 402.710 ;
    END
  END w0_mask_in[291]
  PIN w0_mask_in[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 403.770 0.800 404.070 ;
    END
  END w0_mask_in[292]
  PIN w0_mask_in[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 405.130 0.800 405.430 ;
    END
  END w0_mask_in[293]
  PIN w0_mask_in[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 406.490 0.800 406.790 ;
    END
  END w0_mask_in[294]
  PIN w0_mask_in[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 407.850 0.800 408.150 ;
    END
  END w0_mask_in[295]
  PIN w0_mask_in[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 409.210 0.800 409.510 ;
    END
  END w0_mask_in[296]
  PIN w0_mask_in[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 410.570 0.800 410.870 ;
    END
  END w0_mask_in[297]
  PIN w0_mask_in[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 411.930 0.800 412.230 ;
    END
  END w0_mask_in[298]
  PIN w0_mask_in[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 413.290 0.800 413.590 ;
    END
  END w0_mask_in[299]
  PIN w0_mask_in[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 414.650 0.800 414.950 ;
    END
  END w0_mask_in[300]
  PIN w0_mask_in[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 416.010 0.800 416.310 ;
    END
  END w0_mask_in[301]
  PIN w0_mask_in[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 417.370 0.800 417.670 ;
    END
  END w0_mask_in[302]
  PIN w0_mask_in[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 418.730 0.800 419.030 ;
    END
  END w0_mask_in[303]
  PIN w0_mask_in[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 420.090 0.800 420.390 ;
    END
  END w0_mask_in[304]
  PIN w0_mask_in[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 421.450 0.800 421.750 ;
    END
  END w0_mask_in[305]
  PIN w0_mask_in[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 422.810 0.800 423.110 ;
    END
  END w0_mask_in[306]
  PIN w0_mask_in[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 424.170 0.800 424.470 ;
    END
  END w0_mask_in[307]
  PIN w0_mask_in[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 425.530 0.800 425.830 ;
    END
  END w0_mask_in[308]
  PIN w0_mask_in[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 426.890 0.800 427.190 ;
    END
  END w0_mask_in[309]
  PIN w0_mask_in[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 428.250 0.800 428.550 ;
    END
  END w0_mask_in[310]
  PIN w0_mask_in[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 429.610 0.800 429.910 ;
    END
  END w0_mask_in[311]
  PIN w0_mask_in[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 430.970 0.800 431.270 ;
    END
  END w0_mask_in[312]
  PIN w0_mask_in[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 432.330 0.800 432.630 ;
    END
  END w0_mask_in[313]
  PIN w0_mask_in[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 433.690 0.800 433.990 ;
    END
  END w0_mask_in[314]
  PIN w0_mask_in[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 435.050 0.800 435.350 ;
    END
  END w0_mask_in[315]
  PIN w0_mask_in[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 436.410 0.800 436.710 ;
    END
  END w0_mask_in[316]
  PIN w0_mask_in[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 437.770 0.800 438.070 ;
    END
  END w0_mask_in[317]
  PIN w0_mask_in[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 439.130 0.800 439.430 ;
    END
  END w0_mask_in[318]
  PIN w0_mask_in[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 440.490 0.800 440.790 ;
    END
  END w0_mask_in[319]
  PIN w0_mask_in[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 441.850 0.800 442.150 ;
    END
  END w0_mask_in[320]
  PIN w0_mask_in[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 443.210 0.800 443.510 ;
    END
  END w0_mask_in[321]
  PIN w0_mask_in[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 444.570 0.800 444.870 ;
    END
  END w0_mask_in[322]
  PIN w0_mask_in[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 445.930 0.800 446.230 ;
    END
  END w0_mask_in[323]
  PIN w0_mask_in[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 447.290 0.800 447.590 ;
    END
  END w0_mask_in[324]
  PIN w0_mask_in[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 448.650 0.800 448.950 ;
    END
  END w0_mask_in[325]
  PIN w0_mask_in[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 450.010 0.800 450.310 ;
    END
  END w0_mask_in[326]
  PIN w0_mask_in[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 451.370 0.800 451.670 ;
    END
  END w0_mask_in[327]
  PIN w0_mask_in[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 452.730 0.800 453.030 ;
    END
  END w0_mask_in[328]
  PIN w0_mask_in[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 454.090 0.800 454.390 ;
    END
  END w0_mask_in[329]
  PIN w0_mask_in[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 455.450 0.800 455.750 ;
    END
  END w0_mask_in[330]
  PIN w0_mask_in[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 456.810 0.800 457.110 ;
    END
  END w0_mask_in[331]
  PIN w0_mask_in[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 458.170 0.800 458.470 ;
    END
  END w0_mask_in[332]
  PIN w0_mask_in[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 459.530 0.800 459.830 ;
    END
  END w0_mask_in[333]
  PIN w0_mask_in[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 460.890 0.800 461.190 ;
    END
  END w0_mask_in[334]
  PIN w0_mask_in[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 462.250 0.800 462.550 ;
    END
  END w0_mask_in[335]
  PIN w0_mask_in[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 463.610 0.800 463.910 ;
    END
  END w0_mask_in[336]
  PIN w0_mask_in[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 464.970 0.800 465.270 ;
    END
  END w0_mask_in[337]
  PIN w0_mask_in[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 466.330 0.800 466.630 ;
    END
  END w0_mask_in[338]
  PIN w0_mask_in[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 467.690 0.800 467.990 ;
    END
  END w0_mask_in[339]
  PIN w0_mask_in[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 469.050 0.800 469.350 ;
    END
  END w0_mask_in[340]
  PIN w0_mask_in[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 470.410 0.800 470.710 ;
    END
  END w0_mask_in[341]
  PIN w0_mask_in[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 471.770 0.800 472.070 ;
    END
  END w0_mask_in[342]
  PIN w0_mask_in[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 473.130 0.800 473.430 ;
    END
  END w0_mask_in[343]
  PIN w0_mask_in[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 474.490 0.800 474.790 ;
    END
  END w0_mask_in[344]
  PIN w0_mask_in[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 475.850 0.800 476.150 ;
    END
  END w0_mask_in[345]
  PIN w0_mask_in[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 477.210 0.800 477.510 ;
    END
  END w0_mask_in[346]
  PIN w0_mask_in[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 478.570 0.800 478.870 ;
    END
  END w0_mask_in[347]
  PIN w0_mask_in[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 479.930 0.800 480.230 ;
    END
  END w0_mask_in[348]
  PIN w0_mask_in[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 481.290 0.800 481.590 ;
    END
  END w0_mask_in[349]
  PIN w0_mask_in[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 482.650 0.800 482.950 ;
    END
  END w0_mask_in[350]
  PIN w0_mask_in[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 484.010 0.800 484.310 ;
    END
  END w0_mask_in[351]
  PIN w0_mask_in[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 485.370 0.800 485.670 ;
    END
  END w0_mask_in[352]
  PIN w0_mask_in[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 486.730 0.800 487.030 ;
    END
  END w0_mask_in[353]
  PIN w0_mask_in[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 488.090 0.800 488.390 ;
    END
  END w0_mask_in[354]
  PIN w0_mask_in[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 489.450 0.800 489.750 ;
    END
  END w0_mask_in[355]
  PIN w0_mask_in[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 490.810 0.800 491.110 ;
    END
  END w0_mask_in[356]
  PIN w0_mask_in[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 492.170 0.800 492.470 ;
    END
  END w0_mask_in[357]
  PIN w0_mask_in[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 493.530 0.800 493.830 ;
    END
  END w0_mask_in[358]
  PIN w0_mask_in[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 494.890 0.800 495.190 ;
    END
  END w0_mask_in[359]
  PIN w0_mask_in[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 496.250 0.800 496.550 ;
    END
  END w0_mask_in[360]
  PIN w0_mask_in[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 497.610 0.800 497.910 ;
    END
  END w0_mask_in[361]
  PIN w0_mask_in[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 498.970 0.800 499.270 ;
    END
  END w0_mask_in[362]
  PIN w0_mask_in[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 500.330 0.800 500.630 ;
    END
  END w0_mask_in[363]
  PIN w0_mask_in[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 501.690 0.800 501.990 ;
    END
  END w0_mask_in[364]
  PIN w0_mask_in[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 503.050 0.800 503.350 ;
    END
  END w0_mask_in[365]
  PIN w0_mask_in[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 504.410 0.800 504.710 ;
    END
  END w0_mask_in[366]
  PIN w0_mask_in[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 505.770 0.800 506.070 ;
    END
  END w0_mask_in[367]
  PIN w0_mask_in[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 507.130 0.800 507.430 ;
    END
  END w0_mask_in[368]
  PIN w0_mask_in[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 508.490 0.800 508.790 ;
    END
  END w0_mask_in[369]
  PIN w0_mask_in[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 509.850 0.800 510.150 ;
    END
  END w0_mask_in[370]
  PIN w0_mask_in[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 511.210 0.800 511.510 ;
    END
  END w0_mask_in[371]
  PIN w0_mask_in[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 512.570 0.800 512.870 ;
    END
  END w0_mask_in[372]
  PIN w0_mask_in[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 513.930 0.800 514.230 ;
    END
  END w0_mask_in[373]
  PIN w0_mask_in[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 515.290 0.800 515.590 ;
    END
  END w0_mask_in[374]
  PIN w0_mask_in[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 516.650 0.800 516.950 ;
    END
  END w0_mask_in[375]
  PIN w0_mask_in[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 518.010 0.800 518.310 ;
    END
  END w0_mask_in[376]
  PIN w0_mask_in[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 519.370 0.800 519.670 ;
    END
  END w0_mask_in[377]
  PIN w0_mask_in[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 520.730 0.800 521.030 ;
    END
  END w0_mask_in[378]
  PIN w0_mask_in[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 522.090 0.800 522.390 ;
    END
  END w0_mask_in[379]
  PIN w0_mask_in[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 523.450 0.800 523.750 ;
    END
  END w0_mask_in[380]
  PIN w0_mask_in[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 524.810 0.800 525.110 ;
    END
  END w0_mask_in[381]
  PIN w0_mask_in[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 526.170 0.800 526.470 ;
    END
  END w0_mask_in[382]
  PIN w0_mask_in[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 527.530 0.800 527.830 ;
    END
  END w0_mask_in[383]
  PIN w0_mask_in[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 528.890 0.800 529.190 ;
    END
  END w0_mask_in[384]
  PIN w0_mask_in[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 530.250 0.800 530.550 ;
    END
  END w0_mask_in[385]
  PIN w0_mask_in[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 531.610 0.800 531.910 ;
    END
  END w0_mask_in[386]
  PIN w0_mask_in[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 532.970 0.800 533.270 ;
    END
  END w0_mask_in[387]
  PIN w0_mask_in[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 534.330 0.800 534.630 ;
    END
  END w0_mask_in[388]
  PIN w0_mask_in[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 535.690 0.800 535.990 ;
    END
  END w0_mask_in[389]
  PIN w0_mask_in[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 537.050 0.800 537.350 ;
    END
  END w0_mask_in[390]
  PIN w0_mask_in[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 538.410 0.800 538.710 ;
    END
  END w0_mask_in[391]
  PIN w0_mask_in[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 539.770 0.800 540.070 ;
    END
  END w0_mask_in[392]
  PIN w0_mask_in[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 541.130 0.800 541.430 ;
    END
  END w0_mask_in[393]
  PIN w0_mask_in[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 542.490 0.800 542.790 ;
    END
  END w0_mask_in[394]
  PIN w0_mask_in[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 543.850 0.800 544.150 ;
    END
  END w0_mask_in[395]
  PIN w0_mask_in[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 545.210 0.800 545.510 ;
    END
  END w0_mask_in[396]
  PIN w0_mask_in[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 546.570 0.800 546.870 ;
    END
  END w0_mask_in[397]
  PIN w0_mask_in[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 547.930 0.800 548.230 ;
    END
  END w0_mask_in[398]
  PIN w0_mask_in[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 549.290 0.800 549.590 ;
    END
  END w0_mask_in[399]
  PIN w0_mask_in[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 550.650 0.800 550.950 ;
    END
  END w0_mask_in[400]
  PIN w0_mask_in[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 552.010 0.800 552.310 ;
    END
  END w0_mask_in[401]
  PIN w0_mask_in[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 553.370 0.800 553.670 ;
    END
  END w0_mask_in[402]
  PIN w0_mask_in[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 554.730 0.800 555.030 ;
    END
  END w0_mask_in[403]
  PIN w0_mask_in[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 556.090 0.800 556.390 ;
    END
  END w0_mask_in[404]
  PIN w0_mask_in[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 557.450 0.800 557.750 ;
    END
  END w0_mask_in[405]
  PIN w0_mask_in[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 558.810 0.800 559.110 ;
    END
  END w0_mask_in[406]
  PIN w0_mask_in[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 560.170 0.800 560.470 ;
    END
  END w0_mask_in[407]
  PIN w0_mask_in[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 561.530 0.800 561.830 ;
    END
  END w0_mask_in[408]
  PIN w0_mask_in[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 562.890 0.800 563.190 ;
    END
  END w0_mask_in[409]
  PIN w0_mask_in[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 564.250 0.800 564.550 ;
    END
  END w0_mask_in[410]
  PIN w0_mask_in[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 565.610 0.800 565.910 ;
    END
  END w0_mask_in[411]
  PIN w0_mask_in[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 566.970 0.800 567.270 ;
    END
  END w0_mask_in[412]
  PIN w0_mask_in[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 568.330 0.800 568.630 ;
    END
  END w0_mask_in[413]
  PIN w0_mask_in[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 569.690 0.800 569.990 ;
    END
  END w0_mask_in[414]
  PIN w0_mask_in[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 571.050 0.800 571.350 ;
    END
  END w0_mask_in[415]
  PIN w0_mask_in[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 572.410 0.800 572.710 ;
    END
  END w0_mask_in[416]
  PIN w0_mask_in[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 573.770 0.800 574.070 ;
    END
  END w0_mask_in[417]
  PIN w0_mask_in[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 575.130 0.800 575.430 ;
    END
  END w0_mask_in[418]
  PIN w0_mask_in[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 576.490 0.800 576.790 ;
    END
  END w0_mask_in[419]
  PIN w0_mask_in[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 577.850 0.800 578.150 ;
    END
  END w0_mask_in[420]
  PIN w0_mask_in[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 579.210 0.800 579.510 ;
    END
  END w0_mask_in[421]
  PIN w0_mask_in[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 580.570 0.800 580.870 ;
    END
  END w0_mask_in[422]
  PIN w0_mask_in[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 581.930 0.800 582.230 ;
    END
  END w0_mask_in[423]
  PIN w0_mask_in[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 583.290 0.800 583.590 ;
    END
  END w0_mask_in[424]
  PIN w0_mask_in[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 584.650 0.800 584.950 ;
    END
  END w0_mask_in[425]
  PIN w0_mask_in[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 586.010 0.800 586.310 ;
    END
  END w0_mask_in[426]
  PIN w0_mask_in[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 587.370 0.800 587.670 ;
    END
  END w0_mask_in[427]
  PIN w0_mask_in[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 588.730 0.800 589.030 ;
    END
  END w0_mask_in[428]
  PIN w0_mask_in[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 590.090 0.800 590.390 ;
    END
  END w0_mask_in[429]
  PIN w0_mask_in[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 591.450 0.800 591.750 ;
    END
  END w0_mask_in[430]
  PIN w0_mask_in[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 592.810 0.800 593.110 ;
    END
  END w0_mask_in[431]
  PIN w0_mask_in[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 594.170 0.800 594.470 ;
    END
  END w0_mask_in[432]
  PIN w0_mask_in[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 595.530 0.800 595.830 ;
    END
  END w0_mask_in[433]
  PIN w0_mask_in[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 596.890 0.800 597.190 ;
    END
  END w0_mask_in[434]
  PIN w0_mask_in[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 598.250 0.800 598.550 ;
    END
  END w0_mask_in[435]
  PIN w0_mask_in[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 599.610 0.800 599.910 ;
    END
  END w0_mask_in[436]
  PIN w0_mask_in[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 600.970 0.800 601.270 ;
    END
  END w0_mask_in[437]
  PIN w0_mask_in[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 602.330 0.800 602.630 ;
    END
  END w0_mask_in[438]
  PIN w0_mask_in[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 603.690 0.800 603.990 ;
    END
  END w0_mask_in[439]
  PIN w0_mask_in[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 605.050 0.800 605.350 ;
    END
  END w0_mask_in[440]
  PIN w0_mask_in[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 606.410 0.800 606.710 ;
    END
  END w0_mask_in[441]
  PIN w0_mask_in[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 607.770 0.800 608.070 ;
    END
  END w0_mask_in[442]
  PIN w0_mask_in[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 609.130 0.800 609.430 ;
    END
  END w0_mask_in[443]
  PIN w0_mask_in[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 610.490 0.800 610.790 ;
    END
  END w0_mask_in[444]
  PIN w0_mask_in[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 611.850 0.800 612.150 ;
    END
  END w0_mask_in[445]
  PIN w0_mask_in[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 613.210 0.800 613.510 ;
    END
  END w0_mask_in[446]
  PIN w0_mask_in[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 614.570 0.800 614.870 ;
    END
  END w0_mask_in[447]
  PIN w0_mask_in[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 615.930 0.800 616.230 ;
    END
  END w0_mask_in[448]
  PIN w0_mask_in[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 617.290 0.800 617.590 ;
    END
  END w0_mask_in[449]
  PIN w0_mask_in[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 618.650 0.800 618.950 ;
    END
  END w0_mask_in[450]
  PIN w0_mask_in[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 620.010 0.800 620.310 ;
    END
  END w0_mask_in[451]
  PIN w0_mask_in[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 621.370 0.800 621.670 ;
    END
  END w0_mask_in[452]
  PIN w0_mask_in[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 622.730 0.800 623.030 ;
    END
  END w0_mask_in[453]
  PIN w0_mask_in[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 624.090 0.800 624.390 ;
    END
  END w0_mask_in[454]
  PIN w0_mask_in[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 625.450 0.800 625.750 ;
    END
  END w0_mask_in[455]
  PIN w0_mask_in[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 626.810 0.800 627.110 ;
    END
  END w0_mask_in[456]
  PIN w0_mask_in[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 628.170 0.800 628.470 ;
    END
  END w0_mask_in[457]
  PIN w0_mask_in[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 629.530 0.800 629.830 ;
    END
  END w0_mask_in[458]
  PIN w0_mask_in[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 630.890 0.800 631.190 ;
    END
  END w0_mask_in[459]
  PIN w0_mask_in[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 632.250 0.800 632.550 ;
    END
  END w0_mask_in[460]
  PIN w0_mask_in[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 633.610 0.800 633.910 ;
    END
  END w0_mask_in[461]
  PIN w0_mask_in[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 634.970 0.800 635.270 ;
    END
  END w0_mask_in[462]
  PIN w0_mask_in[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 636.330 0.800 636.630 ;
    END
  END w0_mask_in[463]
  PIN w0_mask_in[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 637.690 0.800 637.990 ;
    END
  END w0_mask_in[464]
  PIN w0_mask_in[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 639.050 0.800 639.350 ;
    END
  END w0_mask_in[465]
  PIN w0_mask_in[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 640.410 0.800 640.710 ;
    END
  END w0_mask_in[466]
  PIN w0_mask_in[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 641.770 0.800 642.070 ;
    END
  END w0_mask_in[467]
  PIN w0_mask_in[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 643.130 0.800 643.430 ;
    END
  END w0_mask_in[468]
  PIN w0_mask_in[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 644.490 0.800 644.790 ;
    END
  END w0_mask_in[469]
  PIN w0_mask_in[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 645.850 0.800 646.150 ;
    END
  END w0_mask_in[470]
  PIN w0_mask_in[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 647.210 0.800 647.510 ;
    END
  END w0_mask_in[471]
  PIN w0_mask_in[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 648.570 0.800 648.870 ;
    END
  END w0_mask_in[472]
  PIN w0_mask_in[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 649.930 0.800 650.230 ;
    END
  END w0_mask_in[473]
  PIN w0_mask_in[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 651.290 0.800 651.590 ;
    END
  END w0_mask_in[474]
  PIN w0_mask_in[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 652.650 0.800 652.950 ;
    END
  END w0_mask_in[475]
  PIN w0_mask_in[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 654.010 0.800 654.310 ;
    END
  END w0_mask_in[476]
  PIN w0_mask_in[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 655.370 0.800 655.670 ;
    END
  END w0_mask_in[477]
  PIN w0_mask_in[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 656.730 0.800 657.030 ;
    END
  END w0_mask_in[478]
  PIN w0_mask_in[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 658.090 0.800 658.390 ;
    END
  END w0_mask_in[479]
  PIN w0_mask_in[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 659.450 0.800 659.750 ;
    END
  END w0_mask_in[480]
  PIN w0_mask_in[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 660.810 0.800 661.110 ;
    END
  END w0_mask_in[481]
  PIN w0_mask_in[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 662.170 0.800 662.470 ;
    END
  END w0_mask_in[482]
  PIN w0_mask_in[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 663.530 0.800 663.830 ;
    END
  END w0_mask_in[483]
  PIN w0_mask_in[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 664.890 0.800 665.190 ;
    END
  END w0_mask_in[484]
  PIN w0_mask_in[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 666.250 0.800 666.550 ;
    END
  END w0_mask_in[485]
  PIN w0_mask_in[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 667.610 0.800 667.910 ;
    END
  END w0_mask_in[486]
  PIN w0_mask_in[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 668.970 0.800 669.270 ;
    END
  END w0_mask_in[487]
  PIN w0_mask_in[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 670.330 0.800 670.630 ;
    END
  END w0_mask_in[488]
  PIN w0_mask_in[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 671.690 0.800 671.990 ;
    END
  END w0_mask_in[489]
  PIN w0_mask_in[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 673.050 0.800 673.350 ;
    END
  END w0_mask_in[490]
  PIN w0_mask_in[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 674.410 0.800 674.710 ;
    END
  END w0_mask_in[491]
  PIN w0_mask_in[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 675.770 0.800 676.070 ;
    END
  END w0_mask_in[492]
  PIN w0_mask_in[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 677.130 0.800 677.430 ;
    END
  END w0_mask_in[493]
  PIN w0_mask_in[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 678.490 0.800 678.790 ;
    END
  END w0_mask_in[494]
  PIN w0_mask_in[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 679.850 0.800 680.150 ;
    END
  END w0_mask_in[495]
  PIN w0_mask_in[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 681.210 0.800 681.510 ;
    END
  END w0_mask_in[496]
  PIN w0_mask_in[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 682.570 0.800 682.870 ;
    END
  END w0_mask_in[497]
  PIN w0_mask_in[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 683.930 0.800 684.230 ;
    END
  END w0_mask_in[498]
  PIN w0_mask_in[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 685.290 0.800 685.590 ;
    END
  END w0_mask_in[499]
  PIN w0_mask_in[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 686.650 0.800 686.950 ;
    END
  END w0_mask_in[500]
  PIN w0_mask_in[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 688.010 0.800 688.310 ;
    END
  END w0_mask_in[501]
  PIN w0_mask_in[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 689.370 0.800 689.670 ;
    END
  END w0_mask_in[502]
  PIN w0_mask_in[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 690.730 0.800 691.030 ;
    END
  END w0_mask_in[503]
  PIN w0_mask_in[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 692.090 0.800 692.390 ;
    END
  END w0_mask_in[504]
  PIN w0_mask_in[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 693.450 0.800 693.750 ;
    END
  END w0_mask_in[505]
  PIN w0_mask_in[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 694.810 0.800 695.110 ;
    END
  END w0_mask_in[506]
  PIN w0_mask_in[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 696.170 0.800 696.470 ;
    END
  END w0_mask_in[507]
  PIN w0_mask_in[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 697.530 0.800 697.830 ;
    END
  END w0_mask_in[508]
  PIN w0_mask_in[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 698.890 0.800 699.190 ;
    END
  END w0_mask_in[509]
  PIN w0_mask_in[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 700.250 0.800 700.550 ;
    END
  END w0_mask_in[510]
  PIN w0_mask_in[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 701.610 0.800 701.910 ;
    END
  END w0_mask_in[511]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 716.570 0.800 716.870 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 717.930 0.800 718.230 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 719.290 0.800 719.590 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 720.650 0.800 720.950 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 722.010 0.800 722.310 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 723.370 0.800 723.670 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 724.730 0.800 725.030 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 726.090 0.800 726.390 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 727.450 0.800 727.750 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 728.810 0.800 729.110 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 730.170 0.800 730.470 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 731.530 0.800 731.830 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 732.890 0.800 733.190 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 734.250 0.800 734.550 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 735.610 0.800 735.910 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 736.970 0.800 737.270 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 738.330 0.800 738.630 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 739.690 0.800 739.990 ;
    END
  END w0_wd_in[17]
  PIN w0_wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 741.050 0.800 741.350 ;
    END
  END w0_wd_in[18]
  PIN w0_wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 742.410 0.800 742.710 ;
    END
  END w0_wd_in[19]
  PIN w0_wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 743.770 0.800 744.070 ;
    END
  END w0_wd_in[20]
  PIN w0_wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 745.130 0.800 745.430 ;
    END
  END w0_wd_in[21]
  PIN w0_wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 746.490 0.800 746.790 ;
    END
  END w0_wd_in[22]
  PIN w0_wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 747.850 0.800 748.150 ;
    END
  END w0_wd_in[23]
  PIN w0_wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 749.210 0.800 749.510 ;
    END
  END w0_wd_in[24]
  PIN w0_wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 750.570 0.800 750.870 ;
    END
  END w0_wd_in[25]
  PIN w0_wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 751.930 0.800 752.230 ;
    END
  END w0_wd_in[26]
  PIN w0_wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 753.290 0.800 753.590 ;
    END
  END w0_wd_in[27]
  PIN w0_wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 754.650 0.800 754.950 ;
    END
  END w0_wd_in[28]
  PIN w0_wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 756.010 0.800 756.310 ;
    END
  END w0_wd_in[29]
  PIN w0_wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 757.370 0.800 757.670 ;
    END
  END w0_wd_in[30]
  PIN w0_wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 758.730 0.800 759.030 ;
    END
  END w0_wd_in[31]
  PIN w0_wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 760.090 0.800 760.390 ;
    END
  END w0_wd_in[32]
  PIN w0_wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 761.450 0.800 761.750 ;
    END
  END w0_wd_in[33]
  PIN w0_wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 762.810 0.800 763.110 ;
    END
  END w0_wd_in[34]
  PIN w0_wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 764.170 0.800 764.470 ;
    END
  END w0_wd_in[35]
  PIN w0_wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 765.530 0.800 765.830 ;
    END
  END w0_wd_in[36]
  PIN w0_wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 766.890 0.800 767.190 ;
    END
  END w0_wd_in[37]
  PIN w0_wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 768.250 0.800 768.550 ;
    END
  END w0_wd_in[38]
  PIN w0_wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 769.610 0.800 769.910 ;
    END
  END w0_wd_in[39]
  PIN w0_wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 770.970 0.800 771.270 ;
    END
  END w0_wd_in[40]
  PIN w0_wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 772.330 0.800 772.630 ;
    END
  END w0_wd_in[41]
  PIN w0_wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 773.690 0.800 773.990 ;
    END
  END w0_wd_in[42]
  PIN w0_wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 775.050 0.800 775.350 ;
    END
  END w0_wd_in[43]
  PIN w0_wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 776.410 0.800 776.710 ;
    END
  END w0_wd_in[44]
  PIN w0_wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 777.770 0.800 778.070 ;
    END
  END w0_wd_in[45]
  PIN w0_wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 779.130 0.800 779.430 ;
    END
  END w0_wd_in[46]
  PIN w0_wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 780.490 0.800 780.790 ;
    END
  END w0_wd_in[47]
  PIN w0_wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 781.850 0.800 782.150 ;
    END
  END w0_wd_in[48]
  PIN w0_wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 783.210 0.800 783.510 ;
    END
  END w0_wd_in[49]
  PIN w0_wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 784.570 0.800 784.870 ;
    END
  END w0_wd_in[50]
  PIN w0_wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 785.930 0.800 786.230 ;
    END
  END w0_wd_in[51]
  PIN w0_wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 787.290 0.800 787.590 ;
    END
  END w0_wd_in[52]
  PIN w0_wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 788.650 0.800 788.950 ;
    END
  END w0_wd_in[53]
  PIN w0_wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 790.010 0.800 790.310 ;
    END
  END w0_wd_in[54]
  PIN w0_wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 791.370 0.800 791.670 ;
    END
  END w0_wd_in[55]
  PIN w0_wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 792.730 0.800 793.030 ;
    END
  END w0_wd_in[56]
  PIN w0_wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 794.090 0.800 794.390 ;
    END
  END w0_wd_in[57]
  PIN w0_wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 795.450 0.800 795.750 ;
    END
  END w0_wd_in[58]
  PIN w0_wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 796.810 0.800 797.110 ;
    END
  END w0_wd_in[59]
  PIN w0_wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 798.170 0.800 798.470 ;
    END
  END w0_wd_in[60]
  PIN w0_wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 799.530 0.800 799.830 ;
    END
  END w0_wd_in[61]
  PIN w0_wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 800.890 0.800 801.190 ;
    END
  END w0_wd_in[62]
  PIN w0_wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 802.250 0.800 802.550 ;
    END
  END w0_wd_in[63]
  PIN w0_wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 803.610 0.800 803.910 ;
    END
  END w0_wd_in[64]
  PIN w0_wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 804.970 0.800 805.270 ;
    END
  END w0_wd_in[65]
  PIN w0_wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 806.330 0.800 806.630 ;
    END
  END w0_wd_in[66]
  PIN w0_wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 807.690 0.800 807.990 ;
    END
  END w0_wd_in[67]
  PIN w0_wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 809.050 0.800 809.350 ;
    END
  END w0_wd_in[68]
  PIN w0_wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 810.410 0.800 810.710 ;
    END
  END w0_wd_in[69]
  PIN w0_wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 811.770 0.800 812.070 ;
    END
  END w0_wd_in[70]
  PIN w0_wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 813.130 0.800 813.430 ;
    END
  END w0_wd_in[71]
  PIN w0_wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 814.490 0.800 814.790 ;
    END
  END w0_wd_in[72]
  PIN w0_wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 815.850 0.800 816.150 ;
    END
  END w0_wd_in[73]
  PIN w0_wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 817.210 0.800 817.510 ;
    END
  END w0_wd_in[74]
  PIN w0_wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 818.570 0.800 818.870 ;
    END
  END w0_wd_in[75]
  PIN w0_wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 819.930 0.800 820.230 ;
    END
  END w0_wd_in[76]
  PIN w0_wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 821.290 0.800 821.590 ;
    END
  END w0_wd_in[77]
  PIN w0_wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 822.650 0.800 822.950 ;
    END
  END w0_wd_in[78]
  PIN w0_wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 824.010 0.800 824.310 ;
    END
  END w0_wd_in[79]
  PIN w0_wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 825.370 0.800 825.670 ;
    END
  END w0_wd_in[80]
  PIN w0_wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 826.730 0.800 827.030 ;
    END
  END w0_wd_in[81]
  PIN w0_wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 828.090 0.800 828.390 ;
    END
  END w0_wd_in[82]
  PIN w0_wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 829.450 0.800 829.750 ;
    END
  END w0_wd_in[83]
  PIN w0_wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 830.810 0.800 831.110 ;
    END
  END w0_wd_in[84]
  PIN w0_wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 832.170 0.800 832.470 ;
    END
  END w0_wd_in[85]
  PIN w0_wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 833.530 0.800 833.830 ;
    END
  END w0_wd_in[86]
  PIN w0_wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 834.890 0.800 835.190 ;
    END
  END w0_wd_in[87]
  PIN w0_wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 836.250 0.800 836.550 ;
    END
  END w0_wd_in[88]
  PIN w0_wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 837.610 0.800 837.910 ;
    END
  END w0_wd_in[89]
  PIN w0_wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 838.970 0.800 839.270 ;
    END
  END w0_wd_in[90]
  PIN w0_wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 840.330 0.800 840.630 ;
    END
  END w0_wd_in[91]
  PIN w0_wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 841.690 0.800 841.990 ;
    END
  END w0_wd_in[92]
  PIN w0_wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 843.050 0.800 843.350 ;
    END
  END w0_wd_in[93]
  PIN w0_wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 844.410 0.800 844.710 ;
    END
  END w0_wd_in[94]
  PIN w0_wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 845.770 0.800 846.070 ;
    END
  END w0_wd_in[95]
  PIN w0_wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 847.130 0.800 847.430 ;
    END
  END w0_wd_in[96]
  PIN w0_wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 848.490 0.800 848.790 ;
    END
  END w0_wd_in[97]
  PIN w0_wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 849.850 0.800 850.150 ;
    END
  END w0_wd_in[98]
  PIN w0_wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 851.210 0.800 851.510 ;
    END
  END w0_wd_in[99]
  PIN w0_wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 852.570 0.800 852.870 ;
    END
  END w0_wd_in[100]
  PIN w0_wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 853.930 0.800 854.230 ;
    END
  END w0_wd_in[101]
  PIN w0_wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 855.290 0.800 855.590 ;
    END
  END w0_wd_in[102]
  PIN w0_wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 856.650 0.800 856.950 ;
    END
  END w0_wd_in[103]
  PIN w0_wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 858.010 0.800 858.310 ;
    END
  END w0_wd_in[104]
  PIN w0_wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 859.370 0.800 859.670 ;
    END
  END w0_wd_in[105]
  PIN w0_wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 860.730 0.800 861.030 ;
    END
  END w0_wd_in[106]
  PIN w0_wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 862.090 0.800 862.390 ;
    END
  END w0_wd_in[107]
  PIN w0_wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 863.450 0.800 863.750 ;
    END
  END w0_wd_in[108]
  PIN w0_wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 864.810 0.800 865.110 ;
    END
  END w0_wd_in[109]
  PIN w0_wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 866.170 0.800 866.470 ;
    END
  END w0_wd_in[110]
  PIN w0_wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 867.530 0.800 867.830 ;
    END
  END w0_wd_in[111]
  PIN w0_wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 868.890 0.800 869.190 ;
    END
  END w0_wd_in[112]
  PIN w0_wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 870.250 0.800 870.550 ;
    END
  END w0_wd_in[113]
  PIN w0_wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 871.610 0.800 871.910 ;
    END
  END w0_wd_in[114]
  PIN w0_wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 872.970 0.800 873.270 ;
    END
  END w0_wd_in[115]
  PIN w0_wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 874.330 0.800 874.630 ;
    END
  END w0_wd_in[116]
  PIN w0_wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 875.690 0.800 875.990 ;
    END
  END w0_wd_in[117]
  PIN w0_wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 877.050 0.800 877.350 ;
    END
  END w0_wd_in[118]
  PIN w0_wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 878.410 0.800 878.710 ;
    END
  END w0_wd_in[119]
  PIN w0_wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 879.770 0.800 880.070 ;
    END
  END w0_wd_in[120]
  PIN w0_wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 881.130 0.800 881.430 ;
    END
  END w0_wd_in[121]
  PIN w0_wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 882.490 0.800 882.790 ;
    END
  END w0_wd_in[122]
  PIN w0_wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 883.850 0.800 884.150 ;
    END
  END w0_wd_in[123]
  PIN w0_wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 885.210 0.800 885.510 ;
    END
  END w0_wd_in[124]
  PIN w0_wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 886.570 0.800 886.870 ;
    END
  END w0_wd_in[125]
  PIN w0_wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 887.930 0.800 888.230 ;
    END
  END w0_wd_in[126]
  PIN w0_wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 889.290 0.800 889.590 ;
    END
  END w0_wd_in[127]
  PIN w0_wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 890.650 0.800 890.950 ;
    END
  END w0_wd_in[128]
  PIN w0_wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 892.010 0.800 892.310 ;
    END
  END w0_wd_in[129]
  PIN w0_wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 893.370 0.800 893.670 ;
    END
  END w0_wd_in[130]
  PIN w0_wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 894.730 0.800 895.030 ;
    END
  END w0_wd_in[131]
  PIN w0_wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 896.090 0.800 896.390 ;
    END
  END w0_wd_in[132]
  PIN w0_wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 897.450 0.800 897.750 ;
    END
  END w0_wd_in[133]
  PIN w0_wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 898.810 0.800 899.110 ;
    END
  END w0_wd_in[134]
  PIN w0_wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 900.170 0.800 900.470 ;
    END
  END w0_wd_in[135]
  PIN w0_wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 901.530 0.800 901.830 ;
    END
  END w0_wd_in[136]
  PIN w0_wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 902.890 0.800 903.190 ;
    END
  END w0_wd_in[137]
  PIN w0_wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 904.250 0.800 904.550 ;
    END
  END w0_wd_in[138]
  PIN w0_wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 905.610 0.800 905.910 ;
    END
  END w0_wd_in[139]
  PIN w0_wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 906.970 0.800 907.270 ;
    END
  END w0_wd_in[140]
  PIN w0_wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 908.330 0.800 908.630 ;
    END
  END w0_wd_in[141]
  PIN w0_wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 909.690 0.800 909.990 ;
    END
  END w0_wd_in[142]
  PIN w0_wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 911.050 0.800 911.350 ;
    END
  END w0_wd_in[143]
  PIN w0_wd_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 912.410 0.800 912.710 ;
    END
  END w0_wd_in[144]
  PIN w0_wd_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 913.770 0.800 914.070 ;
    END
  END w0_wd_in[145]
  PIN w0_wd_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 915.130 0.800 915.430 ;
    END
  END w0_wd_in[146]
  PIN w0_wd_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 916.490 0.800 916.790 ;
    END
  END w0_wd_in[147]
  PIN w0_wd_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 917.850 0.800 918.150 ;
    END
  END w0_wd_in[148]
  PIN w0_wd_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 919.210 0.800 919.510 ;
    END
  END w0_wd_in[149]
  PIN w0_wd_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 920.570 0.800 920.870 ;
    END
  END w0_wd_in[150]
  PIN w0_wd_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 921.930 0.800 922.230 ;
    END
  END w0_wd_in[151]
  PIN w0_wd_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 923.290 0.800 923.590 ;
    END
  END w0_wd_in[152]
  PIN w0_wd_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 924.650 0.800 924.950 ;
    END
  END w0_wd_in[153]
  PIN w0_wd_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 926.010 0.800 926.310 ;
    END
  END w0_wd_in[154]
  PIN w0_wd_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 927.370 0.800 927.670 ;
    END
  END w0_wd_in[155]
  PIN w0_wd_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 928.730 0.800 929.030 ;
    END
  END w0_wd_in[156]
  PIN w0_wd_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 930.090 0.800 930.390 ;
    END
  END w0_wd_in[157]
  PIN w0_wd_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 931.450 0.800 931.750 ;
    END
  END w0_wd_in[158]
  PIN w0_wd_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 932.810 0.800 933.110 ;
    END
  END w0_wd_in[159]
  PIN w0_wd_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 934.170 0.800 934.470 ;
    END
  END w0_wd_in[160]
  PIN w0_wd_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 935.530 0.800 935.830 ;
    END
  END w0_wd_in[161]
  PIN w0_wd_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 936.890 0.800 937.190 ;
    END
  END w0_wd_in[162]
  PIN w0_wd_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 938.250 0.800 938.550 ;
    END
  END w0_wd_in[163]
  PIN w0_wd_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 939.610 0.800 939.910 ;
    END
  END w0_wd_in[164]
  PIN w0_wd_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 940.970 0.800 941.270 ;
    END
  END w0_wd_in[165]
  PIN w0_wd_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 942.330 0.800 942.630 ;
    END
  END w0_wd_in[166]
  PIN w0_wd_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 943.690 0.800 943.990 ;
    END
  END w0_wd_in[167]
  PIN w0_wd_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 945.050 0.800 945.350 ;
    END
  END w0_wd_in[168]
  PIN w0_wd_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 946.410 0.800 946.710 ;
    END
  END w0_wd_in[169]
  PIN w0_wd_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 947.770 0.800 948.070 ;
    END
  END w0_wd_in[170]
  PIN w0_wd_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 949.130 0.800 949.430 ;
    END
  END w0_wd_in[171]
  PIN w0_wd_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 950.490 0.800 950.790 ;
    END
  END w0_wd_in[172]
  PIN w0_wd_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 951.850 0.800 952.150 ;
    END
  END w0_wd_in[173]
  PIN w0_wd_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 953.210 0.800 953.510 ;
    END
  END w0_wd_in[174]
  PIN w0_wd_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 954.570 0.800 954.870 ;
    END
  END w0_wd_in[175]
  PIN w0_wd_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 955.930 0.800 956.230 ;
    END
  END w0_wd_in[176]
  PIN w0_wd_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 957.290 0.800 957.590 ;
    END
  END w0_wd_in[177]
  PIN w0_wd_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 958.650 0.800 958.950 ;
    END
  END w0_wd_in[178]
  PIN w0_wd_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 960.010 0.800 960.310 ;
    END
  END w0_wd_in[179]
  PIN w0_wd_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 961.370 0.800 961.670 ;
    END
  END w0_wd_in[180]
  PIN w0_wd_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 962.730 0.800 963.030 ;
    END
  END w0_wd_in[181]
  PIN w0_wd_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 964.090 0.800 964.390 ;
    END
  END w0_wd_in[182]
  PIN w0_wd_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 965.450 0.800 965.750 ;
    END
  END w0_wd_in[183]
  PIN w0_wd_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 966.810 0.800 967.110 ;
    END
  END w0_wd_in[184]
  PIN w0_wd_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 968.170 0.800 968.470 ;
    END
  END w0_wd_in[185]
  PIN w0_wd_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 969.530 0.800 969.830 ;
    END
  END w0_wd_in[186]
  PIN w0_wd_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 970.890 0.800 971.190 ;
    END
  END w0_wd_in[187]
  PIN w0_wd_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 972.250 0.800 972.550 ;
    END
  END w0_wd_in[188]
  PIN w0_wd_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 973.610 0.800 973.910 ;
    END
  END w0_wd_in[189]
  PIN w0_wd_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 974.970 0.800 975.270 ;
    END
  END w0_wd_in[190]
  PIN w0_wd_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 976.330 0.800 976.630 ;
    END
  END w0_wd_in[191]
  PIN w0_wd_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 977.690 0.800 977.990 ;
    END
  END w0_wd_in[192]
  PIN w0_wd_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 979.050 0.800 979.350 ;
    END
  END w0_wd_in[193]
  PIN w0_wd_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 980.410 0.800 980.710 ;
    END
  END w0_wd_in[194]
  PIN w0_wd_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 981.770 0.800 982.070 ;
    END
  END w0_wd_in[195]
  PIN w0_wd_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 983.130 0.800 983.430 ;
    END
  END w0_wd_in[196]
  PIN w0_wd_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 984.490 0.800 984.790 ;
    END
  END w0_wd_in[197]
  PIN w0_wd_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 985.850 0.800 986.150 ;
    END
  END w0_wd_in[198]
  PIN w0_wd_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 987.210 0.800 987.510 ;
    END
  END w0_wd_in[199]
  PIN w0_wd_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 988.570 0.800 988.870 ;
    END
  END w0_wd_in[200]
  PIN w0_wd_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 989.930 0.800 990.230 ;
    END
  END w0_wd_in[201]
  PIN w0_wd_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 991.290 0.800 991.590 ;
    END
  END w0_wd_in[202]
  PIN w0_wd_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 992.650 0.800 992.950 ;
    END
  END w0_wd_in[203]
  PIN w0_wd_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 994.010 0.800 994.310 ;
    END
  END w0_wd_in[204]
  PIN w0_wd_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 995.370 0.800 995.670 ;
    END
  END w0_wd_in[205]
  PIN w0_wd_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 996.730 0.800 997.030 ;
    END
  END w0_wd_in[206]
  PIN w0_wd_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 998.090 0.800 998.390 ;
    END
  END w0_wd_in[207]
  PIN w0_wd_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 999.450 0.800 999.750 ;
    END
  END w0_wd_in[208]
  PIN w0_wd_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1000.810 0.800 1001.110 ;
    END
  END w0_wd_in[209]
  PIN w0_wd_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1002.170 0.800 1002.470 ;
    END
  END w0_wd_in[210]
  PIN w0_wd_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1003.530 0.800 1003.830 ;
    END
  END w0_wd_in[211]
  PIN w0_wd_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1004.890 0.800 1005.190 ;
    END
  END w0_wd_in[212]
  PIN w0_wd_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1006.250 0.800 1006.550 ;
    END
  END w0_wd_in[213]
  PIN w0_wd_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1007.610 0.800 1007.910 ;
    END
  END w0_wd_in[214]
  PIN w0_wd_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1008.970 0.800 1009.270 ;
    END
  END w0_wd_in[215]
  PIN w0_wd_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1010.330 0.800 1010.630 ;
    END
  END w0_wd_in[216]
  PIN w0_wd_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1011.690 0.800 1011.990 ;
    END
  END w0_wd_in[217]
  PIN w0_wd_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1013.050 0.800 1013.350 ;
    END
  END w0_wd_in[218]
  PIN w0_wd_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1014.410 0.800 1014.710 ;
    END
  END w0_wd_in[219]
  PIN w0_wd_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1015.770 0.800 1016.070 ;
    END
  END w0_wd_in[220]
  PIN w0_wd_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1017.130 0.800 1017.430 ;
    END
  END w0_wd_in[221]
  PIN w0_wd_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1018.490 0.800 1018.790 ;
    END
  END w0_wd_in[222]
  PIN w0_wd_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1019.850 0.800 1020.150 ;
    END
  END w0_wd_in[223]
  PIN w0_wd_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1021.210 0.800 1021.510 ;
    END
  END w0_wd_in[224]
  PIN w0_wd_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1022.570 0.800 1022.870 ;
    END
  END w0_wd_in[225]
  PIN w0_wd_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1023.930 0.800 1024.230 ;
    END
  END w0_wd_in[226]
  PIN w0_wd_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1025.290 0.800 1025.590 ;
    END
  END w0_wd_in[227]
  PIN w0_wd_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1026.650 0.800 1026.950 ;
    END
  END w0_wd_in[228]
  PIN w0_wd_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1028.010 0.800 1028.310 ;
    END
  END w0_wd_in[229]
  PIN w0_wd_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1029.370 0.800 1029.670 ;
    END
  END w0_wd_in[230]
  PIN w0_wd_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1030.730 0.800 1031.030 ;
    END
  END w0_wd_in[231]
  PIN w0_wd_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1032.090 0.800 1032.390 ;
    END
  END w0_wd_in[232]
  PIN w0_wd_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1033.450 0.800 1033.750 ;
    END
  END w0_wd_in[233]
  PIN w0_wd_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1034.810 0.800 1035.110 ;
    END
  END w0_wd_in[234]
  PIN w0_wd_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1036.170 0.800 1036.470 ;
    END
  END w0_wd_in[235]
  PIN w0_wd_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1037.530 0.800 1037.830 ;
    END
  END w0_wd_in[236]
  PIN w0_wd_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1038.890 0.800 1039.190 ;
    END
  END w0_wd_in[237]
  PIN w0_wd_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1040.250 0.800 1040.550 ;
    END
  END w0_wd_in[238]
  PIN w0_wd_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1041.610 0.800 1041.910 ;
    END
  END w0_wd_in[239]
  PIN w0_wd_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1042.970 0.800 1043.270 ;
    END
  END w0_wd_in[240]
  PIN w0_wd_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1044.330 0.800 1044.630 ;
    END
  END w0_wd_in[241]
  PIN w0_wd_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1045.690 0.800 1045.990 ;
    END
  END w0_wd_in[242]
  PIN w0_wd_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1047.050 0.800 1047.350 ;
    END
  END w0_wd_in[243]
  PIN w0_wd_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1048.410 0.800 1048.710 ;
    END
  END w0_wd_in[244]
  PIN w0_wd_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1049.770 0.800 1050.070 ;
    END
  END w0_wd_in[245]
  PIN w0_wd_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1051.130 0.800 1051.430 ;
    END
  END w0_wd_in[246]
  PIN w0_wd_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1052.490 0.800 1052.790 ;
    END
  END w0_wd_in[247]
  PIN w0_wd_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1053.850 0.800 1054.150 ;
    END
  END w0_wd_in[248]
  PIN w0_wd_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1055.210 0.800 1055.510 ;
    END
  END w0_wd_in[249]
  PIN w0_wd_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1056.570 0.800 1056.870 ;
    END
  END w0_wd_in[250]
  PIN w0_wd_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1057.930 0.800 1058.230 ;
    END
  END w0_wd_in[251]
  PIN w0_wd_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1059.290 0.800 1059.590 ;
    END
  END w0_wd_in[252]
  PIN w0_wd_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1060.650 0.800 1060.950 ;
    END
  END w0_wd_in[253]
  PIN w0_wd_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1062.010 0.800 1062.310 ;
    END
  END w0_wd_in[254]
  PIN w0_wd_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1063.370 0.800 1063.670 ;
    END
  END w0_wd_in[255]
  PIN w0_wd_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1064.730 0.800 1065.030 ;
    END
  END w0_wd_in[256]
  PIN w0_wd_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1066.090 0.800 1066.390 ;
    END
  END w0_wd_in[257]
  PIN w0_wd_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1067.450 0.800 1067.750 ;
    END
  END w0_wd_in[258]
  PIN w0_wd_in[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1068.810 0.800 1069.110 ;
    END
  END w0_wd_in[259]
  PIN w0_wd_in[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1070.170 0.800 1070.470 ;
    END
  END w0_wd_in[260]
  PIN w0_wd_in[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1071.530 0.800 1071.830 ;
    END
  END w0_wd_in[261]
  PIN w0_wd_in[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1072.890 0.800 1073.190 ;
    END
  END w0_wd_in[262]
  PIN w0_wd_in[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1074.250 0.800 1074.550 ;
    END
  END w0_wd_in[263]
  PIN w0_wd_in[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1075.610 0.800 1075.910 ;
    END
  END w0_wd_in[264]
  PIN w0_wd_in[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1076.970 0.800 1077.270 ;
    END
  END w0_wd_in[265]
  PIN w0_wd_in[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1078.330 0.800 1078.630 ;
    END
  END w0_wd_in[266]
  PIN w0_wd_in[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1079.690 0.800 1079.990 ;
    END
  END w0_wd_in[267]
  PIN w0_wd_in[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1081.050 0.800 1081.350 ;
    END
  END w0_wd_in[268]
  PIN w0_wd_in[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1082.410 0.800 1082.710 ;
    END
  END w0_wd_in[269]
  PIN w0_wd_in[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1083.770 0.800 1084.070 ;
    END
  END w0_wd_in[270]
  PIN w0_wd_in[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1085.130 0.800 1085.430 ;
    END
  END w0_wd_in[271]
  PIN w0_wd_in[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1086.490 0.800 1086.790 ;
    END
  END w0_wd_in[272]
  PIN w0_wd_in[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1087.850 0.800 1088.150 ;
    END
  END w0_wd_in[273]
  PIN w0_wd_in[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1089.210 0.800 1089.510 ;
    END
  END w0_wd_in[274]
  PIN w0_wd_in[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1090.570 0.800 1090.870 ;
    END
  END w0_wd_in[275]
  PIN w0_wd_in[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1091.930 0.800 1092.230 ;
    END
  END w0_wd_in[276]
  PIN w0_wd_in[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1093.290 0.800 1093.590 ;
    END
  END w0_wd_in[277]
  PIN w0_wd_in[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1094.650 0.800 1094.950 ;
    END
  END w0_wd_in[278]
  PIN w0_wd_in[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1096.010 0.800 1096.310 ;
    END
  END w0_wd_in[279]
  PIN w0_wd_in[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1097.370 0.800 1097.670 ;
    END
  END w0_wd_in[280]
  PIN w0_wd_in[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1098.730 0.800 1099.030 ;
    END
  END w0_wd_in[281]
  PIN w0_wd_in[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1100.090 0.800 1100.390 ;
    END
  END w0_wd_in[282]
  PIN w0_wd_in[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1101.450 0.800 1101.750 ;
    END
  END w0_wd_in[283]
  PIN w0_wd_in[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1102.810 0.800 1103.110 ;
    END
  END w0_wd_in[284]
  PIN w0_wd_in[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1104.170 0.800 1104.470 ;
    END
  END w0_wd_in[285]
  PIN w0_wd_in[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1105.530 0.800 1105.830 ;
    END
  END w0_wd_in[286]
  PIN w0_wd_in[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1106.890 0.800 1107.190 ;
    END
  END w0_wd_in[287]
  PIN w0_wd_in[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1108.250 0.800 1108.550 ;
    END
  END w0_wd_in[288]
  PIN w0_wd_in[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1109.610 0.800 1109.910 ;
    END
  END w0_wd_in[289]
  PIN w0_wd_in[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1110.970 0.800 1111.270 ;
    END
  END w0_wd_in[290]
  PIN w0_wd_in[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1112.330 0.800 1112.630 ;
    END
  END w0_wd_in[291]
  PIN w0_wd_in[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1113.690 0.800 1113.990 ;
    END
  END w0_wd_in[292]
  PIN w0_wd_in[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1115.050 0.800 1115.350 ;
    END
  END w0_wd_in[293]
  PIN w0_wd_in[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1116.410 0.800 1116.710 ;
    END
  END w0_wd_in[294]
  PIN w0_wd_in[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1117.770 0.800 1118.070 ;
    END
  END w0_wd_in[295]
  PIN w0_wd_in[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1119.130 0.800 1119.430 ;
    END
  END w0_wd_in[296]
  PIN w0_wd_in[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1120.490 0.800 1120.790 ;
    END
  END w0_wd_in[297]
  PIN w0_wd_in[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1121.850 0.800 1122.150 ;
    END
  END w0_wd_in[298]
  PIN w0_wd_in[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1123.210 0.800 1123.510 ;
    END
  END w0_wd_in[299]
  PIN w0_wd_in[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1124.570 0.800 1124.870 ;
    END
  END w0_wd_in[300]
  PIN w0_wd_in[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1125.930 0.800 1126.230 ;
    END
  END w0_wd_in[301]
  PIN w0_wd_in[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1127.290 0.800 1127.590 ;
    END
  END w0_wd_in[302]
  PIN w0_wd_in[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1128.650 0.800 1128.950 ;
    END
  END w0_wd_in[303]
  PIN w0_wd_in[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1130.010 0.800 1130.310 ;
    END
  END w0_wd_in[304]
  PIN w0_wd_in[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1131.370 0.800 1131.670 ;
    END
  END w0_wd_in[305]
  PIN w0_wd_in[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1132.730 0.800 1133.030 ;
    END
  END w0_wd_in[306]
  PIN w0_wd_in[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1134.090 0.800 1134.390 ;
    END
  END w0_wd_in[307]
  PIN w0_wd_in[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1135.450 0.800 1135.750 ;
    END
  END w0_wd_in[308]
  PIN w0_wd_in[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1136.810 0.800 1137.110 ;
    END
  END w0_wd_in[309]
  PIN w0_wd_in[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1138.170 0.800 1138.470 ;
    END
  END w0_wd_in[310]
  PIN w0_wd_in[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1139.530 0.800 1139.830 ;
    END
  END w0_wd_in[311]
  PIN w0_wd_in[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1140.890 0.800 1141.190 ;
    END
  END w0_wd_in[312]
  PIN w0_wd_in[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1142.250 0.800 1142.550 ;
    END
  END w0_wd_in[313]
  PIN w0_wd_in[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1143.610 0.800 1143.910 ;
    END
  END w0_wd_in[314]
  PIN w0_wd_in[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1144.970 0.800 1145.270 ;
    END
  END w0_wd_in[315]
  PIN w0_wd_in[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1146.330 0.800 1146.630 ;
    END
  END w0_wd_in[316]
  PIN w0_wd_in[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1147.690 0.800 1147.990 ;
    END
  END w0_wd_in[317]
  PIN w0_wd_in[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1149.050 0.800 1149.350 ;
    END
  END w0_wd_in[318]
  PIN w0_wd_in[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1150.410 0.800 1150.710 ;
    END
  END w0_wd_in[319]
  PIN w0_wd_in[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1151.770 0.800 1152.070 ;
    END
  END w0_wd_in[320]
  PIN w0_wd_in[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1153.130 0.800 1153.430 ;
    END
  END w0_wd_in[321]
  PIN w0_wd_in[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1154.490 0.800 1154.790 ;
    END
  END w0_wd_in[322]
  PIN w0_wd_in[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1155.850 0.800 1156.150 ;
    END
  END w0_wd_in[323]
  PIN w0_wd_in[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1157.210 0.800 1157.510 ;
    END
  END w0_wd_in[324]
  PIN w0_wd_in[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1158.570 0.800 1158.870 ;
    END
  END w0_wd_in[325]
  PIN w0_wd_in[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1159.930 0.800 1160.230 ;
    END
  END w0_wd_in[326]
  PIN w0_wd_in[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1161.290 0.800 1161.590 ;
    END
  END w0_wd_in[327]
  PIN w0_wd_in[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1162.650 0.800 1162.950 ;
    END
  END w0_wd_in[328]
  PIN w0_wd_in[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1164.010 0.800 1164.310 ;
    END
  END w0_wd_in[329]
  PIN w0_wd_in[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1165.370 0.800 1165.670 ;
    END
  END w0_wd_in[330]
  PIN w0_wd_in[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1166.730 0.800 1167.030 ;
    END
  END w0_wd_in[331]
  PIN w0_wd_in[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1168.090 0.800 1168.390 ;
    END
  END w0_wd_in[332]
  PIN w0_wd_in[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1169.450 0.800 1169.750 ;
    END
  END w0_wd_in[333]
  PIN w0_wd_in[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1170.810 0.800 1171.110 ;
    END
  END w0_wd_in[334]
  PIN w0_wd_in[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1172.170 0.800 1172.470 ;
    END
  END w0_wd_in[335]
  PIN w0_wd_in[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1173.530 0.800 1173.830 ;
    END
  END w0_wd_in[336]
  PIN w0_wd_in[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1174.890 0.800 1175.190 ;
    END
  END w0_wd_in[337]
  PIN w0_wd_in[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1176.250 0.800 1176.550 ;
    END
  END w0_wd_in[338]
  PIN w0_wd_in[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1177.610 0.800 1177.910 ;
    END
  END w0_wd_in[339]
  PIN w0_wd_in[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1178.970 0.800 1179.270 ;
    END
  END w0_wd_in[340]
  PIN w0_wd_in[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1180.330 0.800 1180.630 ;
    END
  END w0_wd_in[341]
  PIN w0_wd_in[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1181.690 0.800 1181.990 ;
    END
  END w0_wd_in[342]
  PIN w0_wd_in[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1183.050 0.800 1183.350 ;
    END
  END w0_wd_in[343]
  PIN w0_wd_in[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1184.410 0.800 1184.710 ;
    END
  END w0_wd_in[344]
  PIN w0_wd_in[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1185.770 0.800 1186.070 ;
    END
  END w0_wd_in[345]
  PIN w0_wd_in[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1187.130 0.800 1187.430 ;
    END
  END w0_wd_in[346]
  PIN w0_wd_in[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1188.490 0.800 1188.790 ;
    END
  END w0_wd_in[347]
  PIN w0_wd_in[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1189.850 0.800 1190.150 ;
    END
  END w0_wd_in[348]
  PIN w0_wd_in[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1191.210 0.800 1191.510 ;
    END
  END w0_wd_in[349]
  PIN w0_wd_in[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1192.570 0.800 1192.870 ;
    END
  END w0_wd_in[350]
  PIN w0_wd_in[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1193.930 0.800 1194.230 ;
    END
  END w0_wd_in[351]
  PIN w0_wd_in[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1195.290 0.800 1195.590 ;
    END
  END w0_wd_in[352]
  PIN w0_wd_in[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1196.650 0.800 1196.950 ;
    END
  END w0_wd_in[353]
  PIN w0_wd_in[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1198.010 0.800 1198.310 ;
    END
  END w0_wd_in[354]
  PIN w0_wd_in[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1199.370 0.800 1199.670 ;
    END
  END w0_wd_in[355]
  PIN w0_wd_in[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1200.730 0.800 1201.030 ;
    END
  END w0_wd_in[356]
  PIN w0_wd_in[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1202.090 0.800 1202.390 ;
    END
  END w0_wd_in[357]
  PIN w0_wd_in[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1203.450 0.800 1203.750 ;
    END
  END w0_wd_in[358]
  PIN w0_wd_in[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1204.810 0.800 1205.110 ;
    END
  END w0_wd_in[359]
  PIN w0_wd_in[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1206.170 0.800 1206.470 ;
    END
  END w0_wd_in[360]
  PIN w0_wd_in[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1207.530 0.800 1207.830 ;
    END
  END w0_wd_in[361]
  PIN w0_wd_in[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1208.890 0.800 1209.190 ;
    END
  END w0_wd_in[362]
  PIN w0_wd_in[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1210.250 0.800 1210.550 ;
    END
  END w0_wd_in[363]
  PIN w0_wd_in[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1211.610 0.800 1211.910 ;
    END
  END w0_wd_in[364]
  PIN w0_wd_in[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1212.970 0.800 1213.270 ;
    END
  END w0_wd_in[365]
  PIN w0_wd_in[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1214.330 0.800 1214.630 ;
    END
  END w0_wd_in[366]
  PIN w0_wd_in[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1215.690 0.800 1215.990 ;
    END
  END w0_wd_in[367]
  PIN w0_wd_in[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1217.050 0.800 1217.350 ;
    END
  END w0_wd_in[368]
  PIN w0_wd_in[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1218.410 0.800 1218.710 ;
    END
  END w0_wd_in[369]
  PIN w0_wd_in[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1219.770 0.800 1220.070 ;
    END
  END w0_wd_in[370]
  PIN w0_wd_in[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1221.130 0.800 1221.430 ;
    END
  END w0_wd_in[371]
  PIN w0_wd_in[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1222.490 0.800 1222.790 ;
    END
  END w0_wd_in[372]
  PIN w0_wd_in[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1223.850 0.800 1224.150 ;
    END
  END w0_wd_in[373]
  PIN w0_wd_in[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1225.210 0.800 1225.510 ;
    END
  END w0_wd_in[374]
  PIN w0_wd_in[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1226.570 0.800 1226.870 ;
    END
  END w0_wd_in[375]
  PIN w0_wd_in[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1227.930 0.800 1228.230 ;
    END
  END w0_wd_in[376]
  PIN w0_wd_in[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1229.290 0.800 1229.590 ;
    END
  END w0_wd_in[377]
  PIN w0_wd_in[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1230.650 0.800 1230.950 ;
    END
  END w0_wd_in[378]
  PIN w0_wd_in[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1232.010 0.800 1232.310 ;
    END
  END w0_wd_in[379]
  PIN w0_wd_in[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1233.370 0.800 1233.670 ;
    END
  END w0_wd_in[380]
  PIN w0_wd_in[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1234.730 0.800 1235.030 ;
    END
  END w0_wd_in[381]
  PIN w0_wd_in[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1236.090 0.800 1236.390 ;
    END
  END w0_wd_in[382]
  PIN w0_wd_in[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1237.450 0.800 1237.750 ;
    END
  END w0_wd_in[383]
  PIN w0_wd_in[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1238.810 0.800 1239.110 ;
    END
  END w0_wd_in[384]
  PIN w0_wd_in[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1240.170 0.800 1240.470 ;
    END
  END w0_wd_in[385]
  PIN w0_wd_in[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1241.530 0.800 1241.830 ;
    END
  END w0_wd_in[386]
  PIN w0_wd_in[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1242.890 0.800 1243.190 ;
    END
  END w0_wd_in[387]
  PIN w0_wd_in[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1244.250 0.800 1244.550 ;
    END
  END w0_wd_in[388]
  PIN w0_wd_in[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1245.610 0.800 1245.910 ;
    END
  END w0_wd_in[389]
  PIN w0_wd_in[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1246.970 0.800 1247.270 ;
    END
  END w0_wd_in[390]
  PIN w0_wd_in[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1248.330 0.800 1248.630 ;
    END
  END w0_wd_in[391]
  PIN w0_wd_in[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1249.690 0.800 1249.990 ;
    END
  END w0_wd_in[392]
  PIN w0_wd_in[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1251.050 0.800 1251.350 ;
    END
  END w0_wd_in[393]
  PIN w0_wd_in[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1252.410 0.800 1252.710 ;
    END
  END w0_wd_in[394]
  PIN w0_wd_in[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1253.770 0.800 1254.070 ;
    END
  END w0_wd_in[395]
  PIN w0_wd_in[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1255.130 0.800 1255.430 ;
    END
  END w0_wd_in[396]
  PIN w0_wd_in[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1256.490 0.800 1256.790 ;
    END
  END w0_wd_in[397]
  PIN w0_wd_in[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1257.850 0.800 1258.150 ;
    END
  END w0_wd_in[398]
  PIN w0_wd_in[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1259.210 0.800 1259.510 ;
    END
  END w0_wd_in[399]
  PIN w0_wd_in[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1260.570 0.800 1260.870 ;
    END
  END w0_wd_in[400]
  PIN w0_wd_in[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1261.930 0.800 1262.230 ;
    END
  END w0_wd_in[401]
  PIN w0_wd_in[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1263.290 0.800 1263.590 ;
    END
  END w0_wd_in[402]
  PIN w0_wd_in[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1264.650 0.800 1264.950 ;
    END
  END w0_wd_in[403]
  PIN w0_wd_in[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1266.010 0.800 1266.310 ;
    END
  END w0_wd_in[404]
  PIN w0_wd_in[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1267.370 0.800 1267.670 ;
    END
  END w0_wd_in[405]
  PIN w0_wd_in[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1268.730 0.800 1269.030 ;
    END
  END w0_wd_in[406]
  PIN w0_wd_in[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1270.090 0.800 1270.390 ;
    END
  END w0_wd_in[407]
  PIN w0_wd_in[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1271.450 0.800 1271.750 ;
    END
  END w0_wd_in[408]
  PIN w0_wd_in[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1272.810 0.800 1273.110 ;
    END
  END w0_wd_in[409]
  PIN w0_wd_in[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1274.170 0.800 1274.470 ;
    END
  END w0_wd_in[410]
  PIN w0_wd_in[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1275.530 0.800 1275.830 ;
    END
  END w0_wd_in[411]
  PIN w0_wd_in[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1276.890 0.800 1277.190 ;
    END
  END w0_wd_in[412]
  PIN w0_wd_in[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1278.250 0.800 1278.550 ;
    END
  END w0_wd_in[413]
  PIN w0_wd_in[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1279.610 0.800 1279.910 ;
    END
  END w0_wd_in[414]
  PIN w0_wd_in[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1280.970 0.800 1281.270 ;
    END
  END w0_wd_in[415]
  PIN w0_wd_in[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1282.330 0.800 1282.630 ;
    END
  END w0_wd_in[416]
  PIN w0_wd_in[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1283.690 0.800 1283.990 ;
    END
  END w0_wd_in[417]
  PIN w0_wd_in[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1285.050 0.800 1285.350 ;
    END
  END w0_wd_in[418]
  PIN w0_wd_in[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1286.410 0.800 1286.710 ;
    END
  END w0_wd_in[419]
  PIN w0_wd_in[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1287.770 0.800 1288.070 ;
    END
  END w0_wd_in[420]
  PIN w0_wd_in[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1289.130 0.800 1289.430 ;
    END
  END w0_wd_in[421]
  PIN w0_wd_in[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1290.490 0.800 1290.790 ;
    END
  END w0_wd_in[422]
  PIN w0_wd_in[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1291.850 0.800 1292.150 ;
    END
  END w0_wd_in[423]
  PIN w0_wd_in[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1293.210 0.800 1293.510 ;
    END
  END w0_wd_in[424]
  PIN w0_wd_in[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1294.570 0.800 1294.870 ;
    END
  END w0_wd_in[425]
  PIN w0_wd_in[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1295.930 0.800 1296.230 ;
    END
  END w0_wd_in[426]
  PIN w0_wd_in[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1297.290 0.800 1297.590 ;
    END
  END w0_wd_in[427]
  PIN w0_wd_in[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1298.650 0.800 1298.950 ;
    END
  END w0_wd_in[428]
  PIN w0_wd_in[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1300.010 0.800 1300.310 ;
    END
  END w0_wd_in[429]
  PIN w0_wd_in[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1301.370 0.800 1301.670 ;
    END
  END w0_wd_in[430]
  PIN w0_wd_in[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1302.730 0.800 1303.030 ;
    END
  END w0_wd_in[431]
  PIN w0_wd_in[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1304.090 0.800 1304.390 ;
    END
  END w0_wd_in[432]
  PIN w0_wd_in[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1305.450 0.800 1305.750 ;
    END
  END w0_wd_in[433]
  PIN w0_wd_in[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1306.810 0.800 1307.110 ;
    END
  END w0_wd_in[434]
  PIN w0_wd_in[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1308.170 0.800 1308.470 ;
    END
  END w0_wd_in[435]
  PIN w0_wd_in[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1309.530 0.800 1309.830 ;
    END
  END w0_wd_in[436]
  PIN w0_wd_in[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1310.890 0.800 1311.190 ;
    END
  END w0_wd_in[437]
  PIN w0_wd_in[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1312.250 0.800 1312.550 ;
    END
  END w0_wd_in[438]
  PIN w0_wd_in[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1313.610 0.800 1313.910 ;
    END
  END w0_wd_in[439]
  PIN w0_wd_in[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1314.970 0.800 1315.270 ;
    END
  END w0_wd_in[440]
  PIN w0_wd_in[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1316.330 0.800 1316.630 ;
    END
  END w0_wd_in[441]
  PIN w0_wd_in[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1317.690 0.800 1317.990 ;
    END
  END w0_wd_in[442]
  PIN w0_wd_in[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1319.050 0.800 1319.350 ;
    END
  END w0_wd_in[443]
  PIN w0_wd_in[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1320.410 0.800 1320.710 ;
    END
  END w0_wd_in[444]
  PIN w0_wd_in[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1321.770 0.800 1322.070 ;
    END
  END w0_wd_in[445]
  PIN w0_wd_in[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1323.130 0.800 1323.430 ;
    END
  END w0_wd_in[446]
  PIN w0_wd_in[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1324.490 0.800 1324.790 ;
    END
  END w0_wd_in[447]
  PIN w0_wd_in[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1325.850 0.800 1326.150 ;
    END
  END w0_wd_in[448]
  PIN w0_wd_in[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1327.210 0.800 1327.510 ;
    END
  END w0_wd_in[449]
  PIN w0_wd_in[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1328.570 0.800 1328.870 ;
    END
  END w0_wd_in[450]
  PIN w0_wd_in[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1329.930 0.800 1330.230 ;
    END
  END w0_wd_in[451]
  PIN w0_wd_in[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1331.290 0.800 1331.590 ;
    END
  END w0_wd_in[452]
  PIN w0_wd_in[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1332.650 0.800 1332.950 ;
    END
  END w0_wd_in[453]
  PIN w0_wd_in[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1334.010 0.800 1334.310 ;
    END
  END w0_wd_in[454]
  PIN w0_wd_in[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1335.370 0.800 1335.670 ;
    END
  END w0_wd_in[455]
  PIN w0_wd_in[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1336.730 0.800 1337.030 ;
    END
  END w0_wd_in[456]
  PIN w0_wd_in[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1338.090 0.800 1338.390 ;
    END
  END w0_wd_in[457]
  PIN w0_wd_in[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1339.450 0.800 1339.750 ;
    END
  END w0_wd_in[458]
  PIN w0_wd_in[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1340.810 0.800 1341.110 ;
    END
  END w0_wd_in[459]
  PIN w0_wd_in[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1342.170 0.800 1342.470 ;
    END
  END w0_wd_in[460]
  PIN w0_wd_in[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1343.530 0.800 1343.830 ;
    END
  END w0_wd_in[461]
  PIN w0_wd_in[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1344.890 0.800 1345.190 ;
    END
  END w0_wd_in[462]
  PIN w0_wd_in[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1346.250 0.800 1346.550 ;
    END
  END w0_wd_in[463]
  PIN w0_wd_in[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1347.610 0.800 1347.910 ;
    END
  END w0_wd_in[464]
  PIN w0_wd_in[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1348.970 0.800 1349.270 ;
    END
  END w0_wd_in[465]
  PIN w0_wd_in[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1350.330 0.800 1350.630 ;
    END
  END w0_wd_in[466]
  PIN w0_wd_in[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1351.690 0.800 1351.990 ;
    END
  END w0_wd_in[467]
  PIN w0_wd_in[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1353.050 0.800 1353.350 ;
    END
  END w0_wd_in[468]
  PIN w0_wd_in[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1354.410 0.800 1354.710 ;
    END
  END w0_wd_in[469]
  PIN w0_wd_in[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1355.770 0.800 1356.070 ;
    END
  END w0_wd_in[470]
  PIN w0_wd_in[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1357.130 0.800 1357.430 ;
    END
  END w0_wd_in[471]
  PIN w0_wd_in[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1358.490 0.800 1358.790 ;
    END
  END w0_wd_in[472]
  PIN w0_wd_in[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1359.850 0.800 1360.150 ;
    END
  END w0_wd_in[473]
  PIN w0_wd_in[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1361.210 0.800 1361.510 ;
    END
  END w0_wd_in[474]
  PIN w0_wd_in[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1362.570 0.800 1362.870 ;
    END
  END w0_wd_in[475]
  PIN w0_wd_in[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1363.930 0.800 1364.230 ;
    END
  END w0_wd_in[476]
  PIN w0_wd_in[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1365.290 0.800 1365.590 ;
    END
  END w0_wd_in[477]
  PIN w0_wd_in[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1366.650 0.800 1366.950 ;
    END
  END w0_wd_in[478]
  PIN w0_wd_in[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1368.010 0.800 1368.310 ;
    END
  END w0_wd_in[479]
  PIN w0_wd_in[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1369.370 0.800 1369.670 ;
    END
  END w0_wd_in[480]
  PIN w0_wd_in[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1370.730 0.800 1371.030 ;
    END
  END w0_wd_in[481]
  PIN w0_wd_in[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1372.090 0.800 1372.390 ;
    END
  END w0_wd_in[482]
  PIN w0_wd_in[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1373.450 0.800 1373.750 ;
    END
  END w0_wd_in[483]
  PIN w0_wd_in[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1374.810 0.800 1375.110 ;
    END
  END w0_wd_in[484]
  PIN w0_wd_in[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1376.170 0.800 1376.470 ;
    END
  END w0_wd_in[485]
  PIN w0_wd_in[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1377.530 0.800 1377.830 ;
    END
  END w0_wd_in[486]
  PIN w0_wd_in[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1378.890 0.800 1379.190 ;
    END
  END w0_wd_in[487]
  PIN w0_wd_in[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1380.250 0.800 1380.550 ;
    END
  END w0_wd_in[488]
  PIN w0_wd_in[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1381.610 0.800 1381.910 ;
    END
  END w0_wd_in[489]
  PIN w0_wd_in[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1382.970 0.800 1383.270 ;
    END
  END w0_wd_in[490]
  PIN w0_wd_in[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1384.330 0.800 1384.630 ;
    END
  END w0_wd_in[491]
  PIN w0_wd_in[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1385.690 0.800 1385.990 ;
    END
  END w0_wd_in[492]
  PIN w0_wd_in[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1387.050 0.800 1387.350 ;
    END
  END w0_wd_in[493]
  PIN w0_wd_in[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1388.410 0.800 1388.710 ;
    END
  END w0_wd_in[494]
  PIN w0_wd_in[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1389.770 0.800 1390.070 ;
    END
  END w0_wd_in[495]
  PIN w0_wd_in[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1391.130 0.800 1391.430 ;
    END
  END w0_wd_in[496]
  PIN w0_wd_in[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1392.490 0.800 1392.790 ;
    END
  END w0_wd_in[497]
  PIN w0_wd_in[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1393.850 0.800 1394.150 ;
    END
  END w0_wd_in[498]
  PIN w0_wd_in[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1395.210 0.800 1395.510 ;
    END
  END w0_wd_in[499]
  PIN w0_wd_in[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1396.570 0.800 1396.870 ;
    END
  END w0_wd_in[500]
  PIN w0_wd_in[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1397.930 0.800 1398.230 ;
    END
  END w0_wd_in[501]
  PIN w0_wd_in[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1399.290 0.800 1399.590 ;
    END
  END w0_wd_in[502]
  PIN w0_wd_in[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1400.650 0.800 1400.950 ;
    END
  END w0_wd_in[503]
  PIN w0_wd_in[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1402.010 0.800 1402.310 ;
    END
  END w0_wd_in[504]
  PIN w0_wd_in[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1403.370 0.800 1403.670 ;
    END
  END w0_wd_in[505]
  PIN w0_wd_in[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1404.730 0.800 1405.030 ;
    END
  END w0_wd_in[506]
  PIN w0_wd_in[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1406.090 0.800 1406.390 ;
    END
  END w0_wd_in[507]
  PIN w0_wd_in[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1407.450 0.800 1407.750 ;
    END
  END w0_wd_in[508]
  PIN w0_wd_in[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1408.810 0.800 1409.110 ;
    END
  END w0_wd_in[509]
  PIN w0_wd_in[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1410.170 0.800 1410.470 ;
    END
  END w0_wd_in[510]
  PIN w0_wd_in[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1411.530 0.800 1411.830 ;
    END
  END w0_wd_in[511]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 0.000 4.670 0.350 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 15.570 0.000 15.710 0.350 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 26.610 0.000 26.750 0.350 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 37.650 0.000 37.790 0.350 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 48.690 0.000 48.830 0.350 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 59.730 0.000 59.870 0.350 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 70.770 0.000 70.910 0.350 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 81.810 0.000 81.950 0.350 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 92.850 0.000 92.990 0.350 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 103.890 0.000 104.030 0.350 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 114.930 0.000 115.070 0.350 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 125.970 0.000 126.110 0.350 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 137.010 0.000 137.150 0.350 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 148.050 0.000 148.190 0.350 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 159.090 0.000 159.230 0.350 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 170.130 0.000 170.270 0.350 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 181.170 0.000 181.310 0.350 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 192.210 0.000 192.350 0.350 ;
    END
  END r0_rd_out[17]
  PIN r0_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 203.250 0.000 203.390 0.350 ;
    END
  END r0_rd_out[18]
  PIN r0_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 214.290 0.000 214.430 0.350 ;
    END
  END r0_rd_out[19]
  PIN r0_rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 225.330 0.000 225.470 0.350 ;
    END
  END r0_rd_out[20]
  PIN r0_rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 236.370 0.000 236.510 0.350 ;
    END
  END r0_rd_out[21]
  PIN r0_rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 247.410 0.000 247.550 0.350 ;
    END
  END r0_rd_out[22]
  PIN r0_rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 258.450 0.000 258.590 0.350 ;
    END
  END r0_rd_out[23]
  PIN r0_rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 269.490 0.000 269.630 0.350 ;
    END
  END r0_rd_out[24]
  PIN r0_rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 280.530 0.000 280.670 0.350 ;
    END
  END r0_rd_out[25]
  PIN r0_rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 291.570 0.000 291.710 0.350 ;
    END
  END r0_rd_out[26]
  PIN r0_rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 302.610 0.000 302.750 0.350 ;
    END
  END r0_rd_out[27]
  PIN r0_rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 313.650 0.000 313.790 0.350 ;
    END
  END r0_rd_out[28]
  PIN r0_rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 324.690 0.000 324.830 0.350 ;
    END
  END r0_rd_out[29]
  PIN r0_rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 335.730 0.000 335.870 0.350 ;
    END
  END r0_rd_out[30]
  PIN r0_rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 346.770 0.000 346.910 0.350 ;
    END
  END r0_rd_out[31]
  PIN r0_rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 357.810 0.000 357.950 0.350 ;
    END
  END r0_rd_out[32]
  PIN r0_rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 368.850 0.000 368.990 0.350 ;
    END
  END r0_rd_out[33]
  PIN r0_rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 379.890 0.000 380.030 0.350 ;
    END
  END r0_rd_out[34]
  PIN r0_rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 390.930 0.000 391.070 0.350 ;
    END
  END r0_rd_out[35]
  PIN r0_rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 401.970 0.000 402.110 0.350 ;
    END
  END r0_rd_out[36]
  PIN r0_rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 413.010 0.000 413.150 0.350 ;
    END
  END r0_rd_out[37]
  PIN r0_rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 424.050 0.000 424.190 0.350 ;
    END
  END r0_rd_out[38]
  PIN r0_rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 435.090 0.000 435.230 0.350 ;
    END
  END r0_rd_out[39]
  PIN r0_rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 446.130 0.000 446.270 0.350 ;
    END
  END r0_rd_out[40]
  PIN r0_rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 457.170 0.000 457.310 0.350 ;
    END
  END r0_rd_out[41]
  PIN r0_rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 468.210 0.000 468.350 0.350 ;
    END
  END r0_rd_out[42]
  PIN r0_rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 479.250 0.000 479.390 0.350 ;
    END
  END r0_rd_out[43]
  PIN r0_rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 490.290 0.000 490.430 0.350 ;
    END
  END r0_rd_out[44]
  PIN r0_rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 501.330 0.000 501.470 0.350 ;
    END
  END r0_rd_out[45]
  PIN r0_rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 512.370 0.000 512.510 0.350 ;
    END
  END r0_rd_out[46]
  PIN r0_rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 523.410 0.000 523.550 0.350 ;
    END
  END r0_rd_out[47]
  PIN r0_rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 534.450 0.000 534.590 0.350 ;
    END
  END r0_rd_out[48]
  PIN r0_rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 545.490 0.000 545.630 0.350 ;
    END
  END r0_rd_out[49]
  PIN r0_rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 556.530 0.000 556.670 0.350 ;
    END
  END r0_rd_out[50]
  PIN r0_rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 567.570 0.000 567.710 0.350 ;
    END
  END r0_rd_out[51]
  PIN r0_rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 578.610 0.000 578.750 0.350 ;
    END
  END r0_rd_out[52]
  PIN r0_rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 589.650 0.000 589.790 0.350 ;
    END
  END r0_rd_out[53]
  PIN r0_rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 600.690 0.000 600.830 0.350 ;
    END
  END r0_rd_out[54]
  PIN r0_rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 611.730 0.000 611.870 0.350 ;
    END
  END r0_rd_out[55]
  PIN r0_rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 622.770 0.000 622.910 0.350 ;
    END
  END r0_rd_out[56]
  PIN r0_rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 633.810 0.000 633.950 0.350 ;
    END
  END r0_rd_out[57]
  PIN r0_rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 644.850 0.000 644.990 0.350 ;
    END
  END r0_rd_out[58]
  PIN r0_rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 655.890 0.000 656.030 0.350 ;
    END
  END r0_rd_out[59]
  PIN r0_rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 666.930 0.000 667.070 0.350 ;
    END
  END r0_rd_out[60]
  PIN r0_rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 677.970 0.000 678.110 0.350 ;
    END
  END r0_rd_out[61]
  PIN r0_rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 689.010 0.000 689.150 0.350 ;
    END
  END r0_rd_out[62]
  PIN r0_rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 700.050 0.000 700.190 0.350 ;
    END
  END r0_rd_out[63]
  PIN r0_rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 711.090 0.000 711.230 0.350 ;
    END
  END r0_rd_out[64]
  PIN r0_rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 722.130 0.000 722.270 0.350 ;
    END
  END r0_rd_out[65]
  PIN r0_rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 733.170 0.000 733.310 0.350 ;
    END
  END r0_rd_out[66]
  PIN r0_rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 744.210 0.000 744.350 0.350 ;
    END
  END r0_rd_out[67]
  PIN r0_rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 755.250 0.000 755.390 0.350 ;
    END
  END r0_rd_out[68]
  PIN r0_rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 766.290 0.000 766.430 0.350 ;
    END
  END r0_rd_out[69]
  PIN r0_rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 777.330 0.000 777.470 0.350 ;
    END
  END r0_rd_out[70]
  PIN r0_rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 788.370 0.000 788.510 0.350 ;
    END
  END r0_rd_out[71]
  PIN r0_rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 799.410 0.000 799.550 0.350 ;
    END
  END r0_rd_out[72]
  PIN r0_rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 810.450 0.000 810.590 0.350 ;
    END
  END r0_rd_out[73]
  PIN r0_rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 821.490 0.000 821.630 0.350 ;
    END
  END r0_rd_out[74]
  PIN r0_rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 832.530 0.000 832.670 0.350 ;
    END
  END r0_rd_out[75]
  PIN r0_rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 843.570 0.000 843.710 0.350 ;
    END
  END r0_rd_out[76]
  PIN r0_rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 854.610 0.000 854.750 0.350 ;
    END
  END r0_rd_out[77]
  PIN r0_rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 865.650 0.000 865.790 0.350 ;
    END
  END r0_rd_out[78]
  PIN r0_rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 876.690 0.000 876.830 0.350 ;
    END
  END r0_rd_out[79]
  PIN r0_rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 887.730 0.000 887.870 0.350 ;
    END
  END r0_rd_out[80]
  PIN r0_rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 898.770 0.000 898.910 0.350 ;
    END
  END r0_rd_out[81]
  PIN r0_rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 909.810 0.000 909.950 0.350 ;
    END
  END r0_rd_out[82]
  PIN r0_rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 920.850 0.000 920.990 0.350 ;
    END
  END r0_rd_out[83]
  PIN r0_rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 931.890 0.000 932.030 0.350 ;
    END
  END r0_rd_out[84]
  PIN r0_rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 942.930 0.000 943.070 0.350 ;
    END
  END r0_rd_out[85]
  PIN r0_rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 953.970 0.000 954.110 0.350 ;
    END
  END r0_rd_out[86]
  PIN r0_rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 965.010 0.000 965.150 0.350 ;
    END
  END r0_rd_out[87]
  PIN r0_rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 976.050 0.000 976.190 0.350 ;
    END
  END r0_rd_out[88]
  PIN r0_rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 987.090 0.000 987.230 0.350 ;
    END
  END r0_rd_out[89]
  PIN r0_rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 998.130 0.000 998.270 0.350 ;
    END
  END r0_rd_out[90]
  PIN r0_rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1009.170 0.000 1009.310 0.350 ;
    END
  END r0_rd_out[91]
  PIN r0_rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1020.210 0.000 1020.350 0.350 ;
    END
  END r0_rd_out[92]
  PIN r0_rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1031.250 0.000 1031.390 0.350 ;
    END
  END r0_rd_out[93]
  PIN r0_rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1042.290 0.000 1042.430 0.350 ;
    END
  END r0_rd_out[94]
  PIN r0_rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1053.330 0.000 1053.470 0.350 ;
    END
  END r0_rd_out[95]
  PIN r0_rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1064.370 0.000 1064.510 0.350 ;
    END
  END r0_rd_out[96]
  PIN r0_rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1075.410 0.000 1075.550 0.350 ;
    END
  END r0_rd_out[97]
  PIN r0_rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1086.450 0.000 1086.590 0.350 ;
    END
  END r0_rd_out[98]
  PIN r0_rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1097.490 0.000 1097.630 0.350 ;
    END
  END r0_rd_out[99]
  PIN r0_rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1108.530 0.000 1108.670 0.350 ;
    END
  END r0_rd_out[100]
  PIN r0_rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1119.570 0.000 1119.710 0.350 ;
    END
  END r0_rd_out[101]
  PIN r0_rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1130.610 0.000 1130.750 0.350 ;
    END
  END r0_rd_out[102]
  PIN r0_rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1141.650 0.000 1141.790 0.350 ;
    END
  END r0_rd_out[103]
  PIN r0_rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1152.690 0.000 1152.830 0.350 ;
    END
  END r0_rd_out[104]
  PIN r0_rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1163.730 0.000 1163.870 0.350 ;
    END
  END r0_rd_out[105]
  PIN r0_rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1174.770 0.000 1174.910 0.350 ;
    END
  END r0_rd_out[106]
  PIN r0_rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1185.810 0.000 1185.950 0.350 ;
    END
  END r0_rd_out[107]
  PIN r0_rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1196.850 0.000 1196.990 0.350 ;
    END
  END r0_rd_out[108]
  PIN r0_rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1207.890 0.000 1208.030 0.350 ;
    END
  END r0_rd_out[109]
  PIN r0_rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1218.930 0.000 1219.070 0.350 ;
    END
  END r0_rd_out[110]
  PIN r0_rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1229.970 0.000 1230.110 0.350 ;
    END
  END r0_rd_out[111]
  PIN r0_rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1241.010 0.000 1241.150 0.350 ;
    END
  END r0_rd_out[112]
  PIN r0_rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1252.050 0.000 1252.190 0.350 ;
    END
  END r0_rd_out[113]
  PIN r0_rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1263.090 0.000 1263.230 0.350 ;
    END
  END r0_rd_out[114]
  PIN r0_rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1274.130 0.000 1274.270 0.350 ;
    END
  END r0_rd_out[115]
  PIN r0_rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1285.170 0.000 1285.310 0.350 ;
    END
  END r0_rd_out[116]
  PIN r0_rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1296.210 0.000 1296.350 0.350 ;
    END
  END r0_rd_out[117]
  PIN r0_rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1307.250 0.000 1307.390 0.350 ;
    END
  END r0_rd_out[118]
  PIN r0_rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1318.290 0.000 1318.430 0.350 ;
    END
  END r0_rd_out[119]
  PIN r0_rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1329.330 0.000 1329.470 0.350 ;
    END
  END r0_rd_out[120]
  PIN r0_rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1340.370 0.000 1340.510 0.350 ;
    END
  END r0_rd_out[121]
  PIN r0_rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1351.410 0.000 1351.550 0.350 ;
    END
  END r0_rd_out[122]
  PIN r0_rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1362.450 0.000 1362.590 0.350 ;
    END
  END r0_rd_out[123]
  PIN r0_rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1373.490 0.000 1373.630 0.350 ;
    END
  END r0_rd_out[124]
  PIN r0_rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1384.530 0.000 1384.670 0.350 ;
    END
  END r0_rd_out[125]
  PIN r0_rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1395.570 0.000 1395.710 0.350 ;
    END
  END r0_rd_out[126]
  PIN r0_rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1406.610 0.000 1406.750 0.350 ;
    END
  END r0_rd_out[127]
  PIN r0_rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1417.650 0.000 1417.790 0.350 ;
    END
  END r0_rd_out[128]
  PIN r0_rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1428.690 0.000 1428.830 0.350 ;
    END
  END r0_rd_out[129]
  PIN r0_rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1439.730 0.000 1439.870 0.350 ;
    END
  END r0_rd_out[130]
  PIN r0_rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1450.770 0.000 1450.910 0.350 ;
    END
  END r0_rd_out[131]
  PIN r0_rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1461.810 0.000 1461.950 0.350 ;
    END
  END r0_rd_out[132]
  PIN r0_rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1472.850 0.000 1472.990 0.350 ;
    END
  END r0_rd_out[133]
  PIN r0_rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1483.890 0.000 1484.030 0.350 ;
    END
  END r0_rd_out[134]
  PIN r0_rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1494.930 0.000 1495.070 0.350 ;
    END
  END r0_rd_out[135]
  PIN r0_rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1505.970 0.000 1506.110 0.350 ;
    END
  END r0_rd_out[136]
  PIN r0_rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1517.010 0.000 1517.150 0.350 ;
    END
  END r0_rd_out[137]
  PIN r0_rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1528.050 0.000 1528.190 0.350 ;
    END
  END r0_rd_out[138]
  PIN r0_rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1539.090 0.000 1539.230 0.350 ;
    END
  END r0_rd_out[139]
  PIN r0_rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1550.130 0.000 1550.270 0.350 ;
    END
  END r0_rd_out[140]
  PIN r0_rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1561.170 0.000 1561.310 0.350 ;
    END
  END r0_rd_out[141]
  PIN r0_rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1572.210 0.000 1572.350 0.350 ;
    END
  END r0_rd_out[142]
  PIN r0_rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1583.250 0.000 1583.390 0.350 ;
    END
  END r0_rd_out[143]
  PIN r0_rd_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1594.290 0.000 1594.430 0.350 ;
    END
  END r0_rd_out[144]
  PIN r0_rd_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1605.330 0.000 1605.470 0.350 ;
    END
  END r0_rd_out[145]
  PIN r0_rd_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1616.370 0.000 1616.510 0.350 ;
    END
  END r0_rd_out[146]
  PIN r0_rd_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1627.410 0.000 1627.550 0.350 ;
    END
  END r0_rd_out[147]
  PIN r0_rd_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1638.450 0.000 1638.590 0.350 ;
    END
  END r0_rd_out[148]
  PIN r0_rd_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1649.490 0.000 1649.630 0.350 ;
    END
  END r0_rd_out[149]
  PIN r0_rd_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1660.530 0.000 1660.670 0.350 ;
    END
  END r0_rd_out[150]
  PIN r0_rd_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1671.570 0.000 1671.710 0.350 ;
    END
  END r0_rd_out[151]
  PIN r0_rd_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1682.610 0.000 1682.750 0.350 ;
    END
  END r0_rd_out[152]
  PIN r0_rd_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1693.650 0.000 1693.790 0.350 ;
    END
  END r0_rd_out[153]
  PIN r0_rd_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1704.690 0.000 1704.830 0.350 ;
    END
  END r0_rd_out[154]
  PIN r0_rd_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1715.730 0.000 1715.870 0.350 ;
    END
  END r0_rd_out[155]
  PIN r0_rd_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1726.770 0.000 1726.910 0.350 ;
    END
  END r0_rd_out[156]
  PIN r0_rd_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1737.810 0.000 1737.950 0.350 ;
    END
  END r0_rd_out[157]
  PIN r0_rd_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1748.850 0.000 1748.990 0.350 ;
    END
  END r0_rd_out[158]
  PIN r0_rd_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1759.890 0.000 1760.030 0.350 ;
    END
  END r0_rd_out[159]
  PIN r0_rd_out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1770.930 0.000 1771.070 0.350 ;
    END
  END r0_rd_out[160]
  PIN r0_rd_out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1781.970 0.000 1782.110 0.350 ;
    END
  END r0_rd_out[161]
  PIN r0_rd_out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1793.010 0.000 1793.150 0.350 ;
    END
  END r0_rd_out[162]
  PIN r0_rd_out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1804.050 0.000 1804.190 0.350 ;
    END
  END r0_rd_out[163]
  PIN r0_rd_out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1815.090 0.000 1815.230 0.350 ;
    END
  END r0_rd_out[164]
  PIN r0_rd_out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1826.130 0.000 1826.270 0.350 ;
    END
  END r0_rd_out[165]
  PIN r0_rd_out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1837.170 0.000 1837.310 0.350 ;
    END
  END r0_rd_out[166]
  PIN r0_rd_out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1848.210 0.000 1848.350 0.350 ;
    END
  END r0_rd_out[167]
  PIN r0_rd_out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1859.250 0.000 1859.390 0.350 ;
    END
  END r0_rd_out[168]
  PIN r0_rd_out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1870.290 0.000 1870.430 0.350 ;
    END
  END r0_rd_out[169]
  PIN r0_rd_out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1881.330 0.000 1881.470 0.350 ;
    END
  END r0_rd_out[170]
  PIN r0_rd_out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1892.370 0.000 1892.510 0.350 ;
    END
  END r0_rd_out[171]
  PIN r0_rd_out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1903.410 0.000 1903.550 0.350 ;
    END
  END r0_rd_out[172]
  PIN r0_rd_out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1914.450 0.000 1914.590 0.350 ;
    END
  END r0_rd_out[173]
  PIN r0_rd_out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1925.490 0.000 1925.630 0.350 ;
    END
  END r0_rd_out[174]
  PIN r0_rd_out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1936.530 0.000 1936.670 0.350 ;
    END
  END r0_rd_out[175]
  PIN r0_rd_out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1947.570 0.000 1947.710 0.350 ;
    END
  END r0_rd_out[176]
  PIN r0_rd_out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1958.610 0.000 1958.750 0.350 ;
    END
  END r0_rd_out[177]
  PIN r0_rd_out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1969.650 0.000 1969.790 0.350 ;
    END
  END r0_rd_out[178]
  PIN r0_rd_out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1980.690 0.000 1980.830 0.350 ;
    END
  END r0_rd_out[179]
  PIN r0_rd_out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1991.730 0.000 1991.870 0.350 ;
    END
  END r0_rd_out[180]
  PIN r0_rd_out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2002.770 0.000 2002.910 0.350 ;
    END
  END r0_rd_out[181]
  PIN r0_rd_out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2013.810 0.000 2013.950 0.350 ;
    END
  END r0_rd_out[182]
  PIN r0_rd_out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2024.850 0.000 2024.990 0.350 ;
    END
  END r0_rd_out[183]
  PIN r0_rd_out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2035.890 0.000 2036.030 0.350 ;
    END
  END r0_rd_out[184]
  PIN r0_rd_out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2046.930 0.000 2047.070 0.350 ;
    END
  END r0_rd_out[185]
  PIN r0_rd_out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2057.970 0.000 2058.110 0.350 ;
    END
  END r0_rd_out[186]
  PIN r0_rd_out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2069.010 0.000 2069.150 0.350 ;
    END
  END r0_rd_out[187]
  PIN r0_rd_out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2080.050 0.000 2080.190 0.350 ;
    END
  END r0_rd_out[188]
  PIN r0_rd_out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2091.090 0.000 2091.230 0.350 ;
    END
  END r0_rd_out[189]
  PIN r0_rd_out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2102.130 0.000 2102.270 0.350 ;
    END
  END r0_rd_out[190]
  PIN r0_rd_out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2113.170 0.000 2113.310 0.350 ;
    END
  END r0_rd_out[191]
  PIN r0_rd_out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2124.210 0.000 2124.350 0.350 ;
    END
  END r0_rd_out[192]
  PIN r0_rd_out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2135.250 0.000 2135.390 0.350 ;
    END
  END r0_rd_out[193]
  PIN r0_rd_out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2146.290 0.000 2146.430 0.350 ;
    END
  END r0_rd_out[194]
  PIN r0_rd_out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2157.330 0.000 2157.470 0.350 ;
    END
  END r0_rd_out[195]
  PIN r0_rd_out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2168.370 0.000 2168.510 0.350 ;
    END
  END r0_rd_out[196]
  PIN r0_rd_out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2179.410 0.000 2179.550 0.350 ;
    END
  END r0_rd_out[197]
  PIN r0_rd_out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2190.450 0.000 2190.590 0.350 ;
    END
  END r0_rd_out[198]
  PIN r0_rd_out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2201.490 0.000 2201.630 0.350 ;
    END
  END r0_rd_out[199]
  PIN r0_rd_out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2212.530 0.000 2212.670 0.350 ;
    END
  END r0_rd_out[200]
  PIN r0_rd_out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2223.570 0.000 2223.710 0.350 ;
    END
  END r0_rd_out[201]
  PIN r0_rd_out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2234.610 0.000 2234.750 0.350 ;
    END
  END r0_rd_out[202]
  PIN r0_rd_out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2245.650 0.000 2245.790 0.350 ;
    END
  END r0_rd_out[203]
  PIN r0_rd_out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2256.690 0.000 2256.830 0.350 ;
    END
  END r0_rd_out[204]
  PIN r0_rd_out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2267.730 0.000 2267.870 0.350 ;
    END
  END r0_rd_out[205]
  PIN r0_rd_out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2278.770 0.000 2278.910 0.350 ;
    END
  END r0_rd_out[206]
  PIN r0_rd_out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2289.810 0.000 2289.950 0.350 ;
    END
  END r0_rd_out[207]
  PIN r0_rd_out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2300.850 0.000 2300.990 0.350 ;
    END
  END r0_rd_out[208]
  PIN r0_rd_out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2311.890 0.000 2312.030 0.350 ;
    END
  END r0_rd_out[209]
  PIN r0_rd_out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2322.930 0.000 2323.070 0.350 ;
    END
  END r0_rd_out[210]
  PIN r0_rd_out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2333.970 0.000 2334.110 0.350 ;
    END
  END r0_rd_out[211]
  PIN r0_rd_out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2345.010 0.000 2345.150 0.350 ;
    END
  END r0_rd_out[212]
  PIN r0_rd_out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2356.050 0.000 2356.190 0.350 ;
    END
  END r0_rd_out[213]
  PIN r0_rd_out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2367.090 0.000 2367.230 0.350 ;
    END
  END r0_rd_out[214]
  PIN r0_rd_out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2378.130 0.000 2378.270 0.350 ;
    END
  END r0_rd_out[215]
  PIN r0_rd_out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2389.170 0.000 2389.310 0.350 ;
    END
  END r0_rd_out[216]
  PIN r0_rd_out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2400.210 0.000 2400.350 0.350 ;
    END
  END r0_rd_out[217]
  PIN r0_rd_out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2411.250 0.000 2411.390 0.350 ;
    END
  END r0_rd_out[218]
  PIN r0_rd_out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2422.290 0.000 2422.430 0.350 ;
    END
  END r0_rd_out[219]
  PIN r0_rd_out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2433.330 0.000 2433.470 0.350 ;
    END
  END r0_rd_out[220]
  PIN r0_rd_out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2444.370 0.000 2444.510 0.350 ;
    END
  END r0_rd_out[221]
  PIN r0_rd_out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2455.410 0.000 2455.550 0.350 ;
    END
  END r0_rd_out[222]
  PIN r0_rd_out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2466.450 0.000 2466.590 0.350 ;
    END
  END r0_rd_out[223]
  PIN r0_rd_out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2477.490 0.000 2477.630 0.350 ;
    END
  END r0_rd_out[224]
  PIN r0_rd_out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2488.530 0.000 2488.670 0.350 ;
    END
  END r0_rd_out[225]
  PIN r0_rd_out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2499.570 0.000 2499.710 0.350 ;
    END
  END r0_rd_out[226]
  PIN r0_rd_out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2510.610 0.000 2510.750 0.350 ;
    END
  END r0_rd_out[227]
  PIN r0_rd_out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2521.650 0.000 2521.790 0.350 ;
    END
  END r0_rd_out[228]
  PIN r0_rd_out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2532.690 0.000 2532.830 0.350 ;
    END
  END r0_rd_out[229]
  PIN r0_rd_out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2543.730 0.000 2543.870 0.350 ;
    END
  END r0_rd_out[230]
  PIN r0_rd_out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2554.770 0.000 2554.910 0.350 ;
    END
  END r0_rd_out[231]
  PIN r0_rd_out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2565.810 0.000 2565.950 0.350 ;
    END
  END r0_rd_out[232]
  PIN r0_rd_out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2576.850 0.000 2576.990 0.350 ;
    END
  END r0_rd_out[233]
  PIN r0_rd_out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2587.890 0.000 2588.030 0.350 ;
    END
  END r0_rd_out[234]
  PIN r0_rd_out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2598.930 0.000 2599.070 0.350 ;
    END
  END r0_rd_out[235]
  PIN r0_rd_out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2609.970 0.000 2610.110 0.350 ;
    END
  END r0_rd_out[236]
  PIN r0_rd_out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2621.010 0.000 2621.150 0.350 ;
    END
  END r0_rd_out[237]
  PIN r0_rd_out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2632.050 0.000 2632.190 0.350 ;
    END
  END r0_rd_out[238]
  PIN r0_rd_out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2643.090 0.000 2643.230 0.350 ;
    END
  END r0_rd_out[239]
  PIN r0_rd_out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2654.130 0.000 2654.270 0.350 ;
    END
  END r0_rd_out[240]
  PIN r0_rd_out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2665.170 0.000 2665.310 0.350 ;
    END
  END r0_rd_out[241]
  PIN r0_rd_out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2676.210 0.000 2676.350 0.350 ;
    END
  END r0_rd_out[242]
  PIN r0_rd_out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2687.250 0.000 2687.390 0.350 ;
    END
  END r0_rd_out[243]
  PIN r0_rd_out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2698.290 0.000 2698.430 0.350 ;
    END
  END r0_rd_out[244]
  PIN r0_rd_out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2709.330 0.000 2709.470 0.350 ;
    END
  END r0_rd_out[245]
  PIN r0_rd_out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2720.370 0.000 2720.510 0.350 ;
    END
  END r0_rd_out[246]
  PIN r0_rd_out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2731.410 0.000 2731.550 0.350 ;
    END
  END r0_rd_out[247]
  PIN r0_rd_out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2742.450 0.000 2742.590 0.350 ;
    END
  END r0_rd_out[248]
  PIN r0_rd_out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2753.490 0.000 2753.630 0.350 ;
    END
  END r0_rd_out[249]
  PIN r0_rd_out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2764.530 0.000 2764.670 0.350 ;
    END
  END r0_rd_out[250]
  PIN r0_rd_out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2775.570 0.000 2775.710 0.350 ;
    END
  END r0_rd_out[251]
  PIN r0_rd_out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2786.610 0.000 2786.750 0.350 ;
    END
  END r0_rd_out[252]
  PIN r0_rd_out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2797.650 0.000 2797.790 0.350 ;
    END
  END r0_rd_out[253]
  PIN r0_rd_out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2808.690 0.000 2808.830 0.350 ;
    END
  END r0_rd_out[254]
  PIN r0_rd_out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2819.730 0.000 2819.870 0.350 ;
    END
  END r0_rd_out[255]
  PIN r0_rd_out[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2830.770 0.000 2830.910 0.350 ;
    END
  END r0_rd_out[256]
  PIN r0_rd_out[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2841.810 0.000 2841.950 0.350 ;
    END
  END r0_rd_out[257]
  PIN r0_rd_out[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2852.850 0.000 2852.990 0.350 ;
    END
  END r0_rd_out[258]
  PIN r0_rd_out[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2863.890 0.000 2864.030 0.350 ;
    END
  END r0_rd_out[259]
  PIN r0_rd_out[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2874.930 0.000 2875.070 0.350 ;
    END
  END r0_rd_out[260]
  PIN r0_rd_out[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2885.970 0.000 2886.110 0.350 ;
    END
  END r0_rd_out[261]
  PIN r0_rd_out[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2897.010 0.000 2897.150 0.350 ;
    END
  END r0_rd_out[262]
  PIN r0_rd_out[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2908.050 0.000 2908.190 0.350 ;
    END
  END r0_rd_out[263]
  PIN r0_rd_out[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2919.090 0.000 2919.230 0.350 ;
    END
  END r0_rd_out[264]
  PIN r0_rd_out[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2930.130 0.000 2930.270 0.350 ;
    END
  END r0_rd_out[265]
  PIN r0_rd_out[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2941.170 0.000 2941.310 0.350 ;
    END
  END r0_rd_out[266]
  PIN r0_rd_out[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2952.210 0.000 2952.350 0.350 ;
    END
  END r0_rd_out[267]
  PIN r0_rd_out[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2963.250 0.000 2963.390 0.350 ;
    END
  END r0_rd_out[268]
  PIN r0_rd_out[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2974.290 0.000 2974.430 0.350 ;
    END
  END r0_rd_out[269]
  PIN r0_rd_out[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2985.330 0.000 2985.470 0.350 ;
    END
  END r0_rd_out[270]
  PIN r0_rd_out[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 2996.370 0.000 2996.510 0.350 ;
    END
  END r0_rd_out[271]
  PIN r0_rd_out[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3007.410 0.000 3007.550 0.350 ;
    END
  END r0_rd_out[272]
  PIN r0_rd_out[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3018.450 0.000 3018.590 0.350 ;
    END
  END r0_rd_out[273]
  PIN r0_rd_out[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3029.490 0.000 3029.630 0.350 ;
    END
  END r0_rd_out[274]
  PIN r0_rd_out[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3040.530 0.000 3040.670 0.350 ;
    END
  END r0_rd_out[275]
  PIN r0_rd_out[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3051.570 0.000 3051.710 0.350 ;
    END
  END r0_rd_out[276]
  PIN r0_rd_out[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3062.610 0.000 3062.750 0.350 ;
    END
  END r0_rd_out[277]
  PIN r0_rd_out[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3073.650 0.000 3073.790 0.350 ;
    END
  END r0_rd_out[278]
  PIN r0_rd_out[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3084.690 0.000 3084.830 0.350 ;
    END
  END r0_rd_out[279]
  PIN r0_rd_out[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3095.730 0.000 3095.870 0.350 ;
    END
  END r0_rd_out[280]
  PIN r0_rd_out[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3106.770 0.000 3106.910 0.350 ;
    END
  END r0_rd_out[281]
  PIN r0_rd_out[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3117.810 0.000 3117.950 0.350 ;
    END
  END r0_rd_out[282]
  PIN r0_rd_out[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3128.850 0.000 3128.990 0.350 ;
    END
  END r0_rd_out[283]
  PIN r0_rd_out[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3139.890 0.000 3140.030 0.350 ;
    END
  END r0_rd_out[284]
  PIN r0_rd_out[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3150.930 0.000 3151.070 0.350 ;
    END
  END r0_rd_out[285]
  PIN r0_rd_out[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3161.970 0.000 3162.110 0.350 ;
    END
  END r0_rd_out[286]
  PIN r0_rd_out[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3173.010 0.000 3173.150 0.350 ;
    END
  END r0_rd_out[287]
  PIN r0_rd_out[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3184.050 0.000 3184.190 0.350 ;
    END
  END r0_rd_out[288]
  PIN r0_rd_out[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3195.090 0.000 3195.230 0.350 ;
    END
  END r0_rd_out[289]
  PIN r0_rd_out[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3206.130 0.000 3206.270 0.350 ;
    END
  END r0_rd_out[290]
  PIN r0_rd_out[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3217.170 0.000 3217.310 0.350 ;
    END
  END r0_rd_out[291]
  PIN r0_rd_out[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3228.210 0.000 3228.350 0.350 ;
    END
  END r0_rd_out[292]
  PIN r0_rd_out[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3239.250 0.000 3239.390 0.350 ;
    END
  END r0_rd_out[293]
  PIN r0_rd_out[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3250.290 0.000 3250.430 0.350 ;
    END
  END r0_rd_out[294]
  PIN r0_rd_out[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3261.330 0.000 3261.470 0.350 ;
    END
  END r0_rd_out[295]
  PIN r0_rd_out[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3272.370 0.000 3272.510 0.350 ;
    END
  END r0_rd_out[296]
  PIN r0_rd_out[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3283.410 0.000 3283.550 0.350 ;
    END
  END r0_rd_out[297]
  PIN r0_rd_out[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3294.450 0.000 3294.590 0.350 ;
    END
  END r0_rd_out[298]
  PIN r0_rd_out[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3305.490 0.000 3305.630 0.350 ;
    END
  END r0_rd_out[299]
  PIN r0_rd_out[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3316.530 0.000 3316.670 0.350 ;
    END
  END r0_rd_out[300]
  PIN r0_rd_out[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3327.570 0.000 3327.710 0.350 ;
    END
  END r0_rd_out[301]
  PIN r0_rd_out[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3338.610 0.000 3338.750 0.350 ;
    END
  END r0_rd_out[302]
  PIN r0_rd_out[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3349.650 0.000 3349.790 0.350 ;
    END
  END r0_rd_out[303]
  PIN r0_rd_out[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3360.690 0.000 3360.830 0.350 ;
    END
  END r0_rd_out[304]
  PIN r0_rd_out[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3371.730 0.000 3371.870 0.350 ;
    END
  END r0_rd_out[305]
  PIN r0_rd_out[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3382.770 0.000 3382.910 0.350 ;
    END
  END r0_rd_out[306]
  PIN r0_rd_out[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3393.810 0.000 3393.950 0.350 ;
    END
  END r0_rd_out[307]
  PIN r0_rd_out[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3404.850 0.000 3404.990 0.350 ;
    END
  END r0_rd_out[308]
  PIN r0_rd_out[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3415.890 0.000 3416.030 0.350 ;
    END
  END r0_rd_out[309]
  PIN r0_rd_out[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3426.930 0.000 3427.070 0.350 ;
    END
  END r0_rd_out[310]
  PIN r0_rd_out[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3437.970 0.000 3438.110 0.350 ;
    END
  END r0_rd_out[311]
  PIN r0_rd_out[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3449.010 0.000 3449.150 0.350 ;
    END
  END r0_rd_out[312]
  PIN r0_rd_out[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3460.050 0.000 3460.190 0.350 ;
    END
  END r0_rd_out[313]
  PIN r0_rd_out[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3471.090 0.000 3471.230 0.350 ;
    END
  END r0_rd_out[314]
  PIN r0_rd_out[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3482.130 0.000 3482.270 0.350 ;
    END
  END r0_rd_out[315]
  PIN r0_rd_out[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3493.170 0.000 3493.310 0.350 ;
    END
  END r0_rd_out[316]
  PIN r0_rd_out[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3504.210 0.000 3504.350 0.350 ;
    END
  END r0_rd_out[317]
  PIN r0_rd_out[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3515.250 0.000 3515.390 0.350 ;
    END
  END r0_rd_out[318]
  PIN r0_rd_out[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3526.290 0.000 3526.430 0.350 ;
    END
  END r0_rd_out[319]
  PIN r0_rd_out[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3537.330 0.000 3537.470 0.350 ;
    END
  END r0_rd_out[320]
  PIN r0_rd_out[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3548.370 0.000 3548.510 0.350 ;
    END
  END r0_rd_out[321]
  PIN r0_rd_out[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3559.410 0.000 3559.550 0.350 ;
    END
  END r0_rd_out[322]
  PIN r0_rd_out[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3570.450 0.000 3570.590 0.350 ;
    END
  END r0_rd_out[323]
  PIN r0_rd_out[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3581.490 0.000 3581.630 0.350 ;
    END
  END r0_rd_out[324]
  PIN r0_rd_out[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3592.530 0.000 3592.670 0.350 ;
    END
  END r0_rd_out[325]
  PIN r0_rd_out[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3603.570 0.000 3603.710 0.350 ;
    END
  END r0_rd_out[326]
  PIN r0_rd_out[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3614.610 0.000 3614.750 0.350 ;
    END
  END r0_rd_out[327]
  PIN r0_rd_out[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3625.650 0.000 3625.790 0.350 ;
    END
  END r0_rd_out[328]
  PIN r0_rd_out[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3636.690 0.000 3636.830 0.350 ;
    END
  END r0_rd_out[329]
  PIN r0_rd_out[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3647.730 0.000 3647.870 0.350 ;
    END
  END r0_rd_out[330]
  PIN r0_rd_out[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3658.770 0.000 3658.910 0.350 ;
    END
  END r0_rd_out[331]
  PIN r0_rd_out[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3669.810 0.000 3669.950 0.350 ;
    END
  END r0_rd_out[332]
  PIN r0_rd_out[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3680.850 0.000 3680.990 0.350 ;
    END
  END r0_rd_out[333]
  PIN r0_rd_out[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3691.890 0.000 3692.030 0.350 ;
    END
  END r0_rd_out[334]
  PIN r0_rd_out[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3702.930 0.000 3703.070 0.350 ;
    END
  END r0_rd_out[335]
  PIN r0_rd_out[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3713.970 0.000 3714.110 0.350 ;
    END
  END r0_rd_out[336]
  PIN r0_rd_out[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3725.010 0.000 3725.150 0.350 ;
    END
  END r0_rd_out[337]
  PIN r0_rd_out[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3736.050 0.000 3736.190 0.350 ;
    END
  END r0_rd_out[338]
  PIN r0_rd_out[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3747.090 0.000 3747.230 0.350 ;
    END
  END r0_rd_out[339]
  PIN r0_rd_out[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3758.130 0.000 3758.270 0.350 ;
    END
  END r0_rd_out[340]
  PIN r0_rd_out[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3769.170 0.000 3769.310 0.350 ;
    END
  END r0_rd_out[341]
  PIN r0_rd_out[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3780.210 0.000 3780.350 0.350 ;
    END
  END r0_rd_out[342]
  PIN r0_rd_out[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3791.250 0.000 3791.390 0.350 ;
    END
  END r0_rd_out[343]
  PIN r0_rd_out[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3802.290 0.000 3802.430 0.350 ;
    END
  END r0_rd_out[344]
  PIN r0_rd_out[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3813.330 0.000 3813.470 0.350 ;
    END
  END r0_rd_out[345]
  PIN r0_rd_out[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3824.370 0.000 3824.510 0.350 ;
    END
  END r0_rd_out[346]
  PIN r0_rd_out[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3835.410 0.000 3835.550 0.350 ;
    END
  END r0_rd_out[347]
  PIN r0_rd_out[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3846.450 0.000 3846.590 0.350 ;
    END
  END r0_rd_out[348]
  PIN r0_rd_out[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3857.490 0.000 3857.630 0.350 ;
    END
  END r0_rd_out[349]
  PIN r0_rd_out[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3868.530 0.000 3868.670 0.350 ;
    END
  END r0_rd_out[350]
  PIN r0_rd_out[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3879.570 0.000 3879.710 0.350 ;
    END
  END r0_rd_out[351]
  PIN r0_rd_out[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3890.610 0.000 3890.750 0.350 ;
    END
  END r0_rd_out[352]
  PIN r0_rd_out[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3901.650 0.000 3901.790 0.350 ;
    END
  END r0_rd_out[353]
  PIN r0_rd_out[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3912.690 0.000 3912.830 0.350 ;
    END
  END r0_rd_out[354]
  PIN r0_rd_out[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3923.730 0.000 3923.870 0.350 ;
    END
  END r0_rd_out[355]
  PIN r0_rd_out[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3934.770 0.000 3934.910 0.350 ;
    END
  END r0_rd_out[356]
  PIN r0_rd_out[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3945.810 0.000 3945.950 0.350 ;
    END
  END r0_rd_out[357]
  PIN r0_rd_out[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3956.850 0.000 3956.990 0.350 ;
    END
  END r0_rd_out[358]
  PIN r0_rd_out[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3967.890 0.000 3968.030 0.350 ;
    END
  END r0_rd_out[359]
  PIN r0_rd_out[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3978.930 0.000 3979.070 0.350 ;
    END
  END r0_rd_out[360]
  PIN r0_rd_out[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 3989.970 0.000 3990.110 0.350 ;
    END
  END r0_rd_out[361]
  PIN r0_rd_out[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4001.010 0.000 4001.150 0.350 ;
    END
  END r0_rd_out[362]
  PIN r0_rd_out[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4012.050 0.000 4012.190 0.350 ;
    END
  END r0_rd_out[363]
  PIN r0_rd_out[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4023.090 0.000 4023.230 0.350 ;
    END
  END r0_rd_out[364]
  PIN r0_rd_out[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4034.130 0.000 4034.270 0.350 ;
    END
  END r0_rd_out[365]
  PIN r0_rd_out[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4045.170 0.000 4045.310 0.350 ;
    END
  END r0_rd_out[366]
  PIN r0_rd_out[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4056.210 0.000 4056.350 0.350 ;
    END
  END r0_rd_out[367]
  PIN r0_rd_out[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4067.250 0.000 4067.390 0.350 ;
    END
  END r0_rd_out[368]
  PIN r0_rd_out[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4078.290 0.000 4078.430 0.350 ;
    END
  END r0_rd_out[369]
  PIN r0_rd_out[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4089.330 0.000 4089.470 0.350 ;
    END
  END r0_rd_out[370]
  PIN r0_rd_out[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4100.370 0.000 4100.510 0.350 ;
    END
  END r0_rd_out[371]
  PIN r0_rd_out[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4111.410 0.000 4111.550 0.350 ;
    END
  END r0_rd_out[372]
  PIN r0_rd_out[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4122.450 0.000 4122.590 0.350 ;
    END
  END r0_rd_out[373]
  PIN r0_rd_out[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4133.490 0.000 4133.630 0.350 ;
    END
  END r0_rd_out[374]
  PIN r0_rd_out[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4144.530 0.000 4144.670 0.350 ;
    END
  END r0_rd_out[375]
  PIN r0_rd_out[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4155.570 0.000 4155.710 0.350 ;
    END
  END r0_rd_out[376]
  PIN r0_rd_out[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4166.610 0.000 4166.750 0.350 ;
    END
  END r0_rd_out[377]
  PIN r0_rd_out[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4177.650 0.000 4177.790 0.350 ;
    END
  END r0_rd_out[378]
  PIN r0_rd_out[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4188.690 0.000 4188.830 0.350 ;
    END
  END r0_rd_out[379]
  PIN r0_rd_out[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4199.730 0.000 4199.870 0.350 ;
    END
  END r0_rd_out[380]
  PIN r0_rd_out[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4210.770 0.000 4210.910 0.350 ;
    END
  END r0_rd_out[381]
  PIN r0_rd_out[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4221.810 0.000 4221.950 0.350 ;
    END
  END r0_rd_out[382]
  PIN r0_rd_out[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4232.850 0.000 4232.990 0.350 ;
    END
  END r0_rd_out[383]
  PIN r0_rd_out[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4243.890 0.000 4244.030 0.350 ;
    END
  END r0_rd_out[384]
  PIN r0_rd_out[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4254.930 0.000 4255.070 0.350 ;
    END
  END r0_rd_out[385]
  PIN r0_rd_out[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4265.970 0.000 4266.110 0.350 ;
    END
  END r0_rd_out[386]
  PIN r0_rd_out[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4277.010 0.000 4277.150 0.350 ;
    END
  END r0_rd_out[387]
  PIN r0_rd_out[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4288.050 0.000 4288.190 0.350 ;
    END
  END r0_rd_out[388]
  PIN r0_rd_out[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4299.090 0.000 4299.230 0.350 ;
    END
  END r0_rd_out[389]
  PIN r0_rd_out[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4310.130 0.000 4310.270 0.350 ;
    END
  END r0_rd_out[390]
  PIN r0_rd_out[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4321.170 0.000 4321.310 0.350 ;
    END
  END r0_rd_out[391]
  PIN r0_rd_out[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4332.210 0.000 4332.350 0.350 ;
    END
  END r0_rd_out[392]
  PIN r0_rd_out[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4343.250 0.000 4343.390 0.350 ;
    END
  END r0_rd_out[393]
  PIN r0_rd_out[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4354.290 0.000 4354.430 0.350 ;
    END
  END r0_rd_out[394]
  PIN r0_rd_out[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4365.330 0.000 4365.470 0.350 ;
    END
  END r0_rd_out[395]
  PIN r0_rd_out[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4376.370 0.000 4376.510 0.350 ;
    END
  END r0_rd_out[396]
  PIN r0_rd_out[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4387.410 0.000 4387.550 0.350 ;
    END
  END r0_rd_out[397]
  PIN r0_rd_out[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4398.450 0.000 4398.590 0.350 ;
    END
  END r0_rd_out[398]
  PIN r0_rd_out[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4409.490 0.000 4409.630 0.350 ;
    END
  END r0_rd_out[399]
  PIN r0_rd_out[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4420.530 0.000 4420.670 0.350 ;
    END
  END r0_rd_out[400]
  PIN r0_rd_out[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4431.570 0.000 4431.710 0.350 ;
    END
  END r0_rd_out[401]
  PIN r0_rd_out[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4442.610 0.000 4442.750 0.350 ;
    END
  END r0_rd_out[402]
  PIN r0_rd_out[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4453.650 0.000 4453.790 0.350 ;
    END
  END r0_rd_out[403]
  PIN r0_rd_out[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4464.690 0.000 4464.830 0.350 ;
    END
  END r0_rd_out[404]
  PIN r0_rd_out[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4475.730 0.000 4475.870 0.350 ;
    END
  END r0_rd_out[405]
  PIN r0_rd_out[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4486.770 0.000 4486.910 0.350 ;
    END
  END r0_rd_out[406]
  PIN r0_rd_out[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4497.810 0.000 4497.950 0.350 ;
    END
  END r0_rd_out[407]
  PIN r0_rd_out[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4508.850 0.000 4508.990 0.350 ;
    END
  END r0_rd_out[408]
  PIN r0_rd_out[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4519.890 0.000 4520.030 0.350 ;
    END
  END r0_rd_out[409]
  PIN r0_rd_out[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4530.930 0.000 4531.070 0.350 ;
    END
  END r0_rd_out[410]
  PIN r0_rd_out[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4541.970 0.000 4542.110 0.350 ;
    END
  END r0_rd_out[411]
  PIN r0_rd_out[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4553.010 0.000 4553.150 0.350 ;
    END
  END r0_rd_out[412]
  PIN r0_rd_out[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4564.050 0.000 4564.190 0.350 ;
    END
  END r0_rd_out[413]
  PIN r0_rd_out[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4575.090 0.000 4575.230 0.350 ;
    END
  END r0_rd_out[414]
  PIN r0_rd_out[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4586.130 0.000 4586.270 0.350 ;
    END
  END r0_rd_out[415]
  PIN r0_rd_out[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4597.170 0.000 4597.310 0.350 ;
    END
  END r0_rd_out[416]
  PIN r0_rd_out[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4608.210 0.000 4608.350 0.350 ;
    END
  END r0_rd_out[417]
  PIN r0_rd_out[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4619.250 0.000 4619.390 0.350 ;
    END
  END r0_rd_out[418]
  PIN r0_rd_out[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4630.290 0.000 4630.430 0.350 ;
    END
  END r0_rd_out[419]
  PIN r0_rd_out[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4641.330 0.000 4641.470 0.350 ;
    END
  END r0_rd_out[420]
  PIN r0_rd_out[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4652.370 0.000 4652.510 0.350 ;
    END
  END r0_rd_out[421]
  PIN r0_rd_out[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4663.410 0.000 4663.550 0.350 ;
    END
  END r0_rd_out[422]
  PIN r0_rd_out[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4674.450 0.000 4674.590 0.350 ;
    END
  END r0_rd_out[423]
  PIN r0_rd_out[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4685.490 0.000 4685.630 0.350 ;
    END
  END r0_rd_out[424]
  PIN r0_rd_out[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4696.530 0.000 4696.670 0.350 ;
    END
  END r0_rd_out[425]
  PIN r0_rd_out[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4707.570 0.000 4707.710 0.350 ;
    END
  END r0_rd_out[426]
  PIN r0_rd_out[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4718.610 0.000 4718.750 0.350 ;
    END
  END r0_rd_out[427]
  PIN r0_rd_out[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4729.650 0.000 4729.790 0.350 ;
    END
  END r0_rd_out[428]
  PIN r0_rd_out[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4740.690 0.000 4740.830 0.350 ;
    END
  END r0_rd_out[429]
  PIN r0_rd_out[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4751.730 0.000 4751.870 0.350 ;
    END
  END r0_rd_out[430]
  PIN r0_rd_out[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4762.770 0.000 4762.910 0.350 ;
    END
  END r0_rd_out[431]
  PIN r0_rd_out[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4773.810 0.000 4773.950 0.350 ;
    END
  END r0_rd_out[432]
  PIN r0_rd_out[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4784.850 0.000 4784.990 0.350 ;
    END
  END r0_rd_out[433]
  PIN r0_rd_out[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4795.890 0.000 4796.030 0.350 ;
    END
  END r0_rd_out[434]
  PIN r0_rd_out[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4806.930 0.000 4807.070 0.350 ;
    END
  END r0_rd_out[435]
  PIN r0_rd_out[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4817.970 0.000 4818.110 0.350 ;
    END
  END r0_rd_out[436]
  PIN r0_rd_out[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4829.010 0.000 4829.150 0.350 ;
    END
  END r0_rd_out[437]
  PIN r0_rd_out[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4840.050 0.000 4840.190 0.350 ;
    END
  END r0_rd_out[438]
  PIN r0_rd_out[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4851.090 0.000 4851.230 0.350 ;
    END
  END r0_rd_out[439]
  PIN r0_rd_out[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4862.130 0.000 4862.270 0.350 ;
    END
  END r0_rd_out[440]
  PIN r0_rd_out[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4873.170 0.000 4873.310 0.350 ;
    END
  END r0_rd_out[441]
  PIN r0_rd_out[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4884.210 0.000 4884.350 0.350 ;
    END
  END r0_rd_out[442]
  PIN r0_rd_out[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4895.250 0.000 4895.390 0.350 ;
    END
  END r0_rd_out[443]
  PIN r0_rd_out[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4906.290 0.000 4906.430 0.350 ;
    END
  END r0_rd_out[444]
  PIN r0_rd_out[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4917.330 0.000 4917.470 0.350 ;
    END
  END r0_rd_out[445]
  PIN r0_rd_out[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4928.370 0.000 4928.510 0.350 ;
    END
  END r0_rd_out[446]
  PIN r0_rd_out[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4939.410 0.000 4939.550 0.350 ;
    END
  END r0_rd_out[447]
  PIN r0_rd_out[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4950.450 0.000 4950.590 0.350 ;
    END
  END r0_rd_out[448]
  PIN r0_rd_out[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4961.490 0.000 4961.630 0.350 ;
    END
  END r0_rd_out[449]
  PIN r0_rd_out[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4972.530 0.000 4972.670 0.350 ;
    END
  END r0_rd_out[450]
  PIN r0_rd_out[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4983.570 0.000 4983.710 0.350 ;
    END
  END r0_rd_out[451]
  PIN r0_rd_out[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4994.610 0.000 4994.750 0.350 ;
    END
  END r0_rd_out[452]
  PIN r0_rd_out[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5005.650 0.000 5005.790 0.350 ;
    END
  END r0_rd_out[453]
  PIN r0_rd_out[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5016.690 0.000 5016.830 0.350 ;
    END
  END r0_rd_out[454]
  PIN r0_rd_out[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5027.730 0.000 5027.870 0.350 ;
    END
  END r0_rd_out[455]
  PIN r0_rd_out[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5038.770 0.000 5038.910 0.350 ;
    END
  END r0_rd_out[456]
  PIN r0_rd_out[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5049.810 0.000 5049.950 0.350 ;
    END
  END r0_rd_out[457]
  PIN r0_rd_out[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5060.850 0.000 5060.990 0.350 ;
    END
  END r0_rd_out[458]
  PIN r0_rd_out[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5071.890 0.000 5072.030 0.350 ;
    END
  END r0_rd_out[459]
  PIN r0_rd_out[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5082.930 0.000 5083.070 0.350 ;
    END
  END r0_rd_out[460]
  PIN r0_rd_out[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5093.970 0.000 5094.110 0.350 ;
    END
  END r0_rd_out[461]
  PIN r0_rd_out[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5105.010 0.000 5105.150 0.350 ;
    END
  END r0_rd_out[462]
  PIN r0_rd_out[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5116.050 0.000 5116.190 0.350 ;
    END
  END r0_rd_out[463]
  PIN r0_rd_out[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5127.090 0.000 5127.230 0.350 ;
    END
  END r0_rd_out[464]
  PIN r0_rd_out[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5138.130 0.000 5138.270 0.350 ;
    END
  END r0_rd_out[465]
  PIN r0_rd_out[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5149.170 0.000 5149.310 0.350 ;
    END
  END r0_rd_out[466]
  PIN r0_rd_out[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5160.210 0.000 5160.350 0.350 ;
    END
  END r0_rd_out[467]
  PIN r0_rd_out[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5171.250 0.000 5171.390 0.350 ;
    END
  END r0_rd_out[468]
  PIN r0_rd_out[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5182.290 0.000 5182.430 0.350 ;
    END
  END r0_rd_out[469]
  PIN r0_rd_out[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5193.330 0.000 5193.470 0.350 ;
    END
  END r0_rd_out[470]
  PIN r0_rd_out[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5204.370 0.000 5204.510 0.350 ;
    END
  END r0_rd_out[471]
  PIN r0_rd_out[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5215.410 0.000 5215.550 0.350 ;
    END
  END r0_rd_out[472]
  PIN r0_rd_out[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5226.450 0.000 5226.590 0.350 ;
    END
  END r0_rd_out[473]
  PIN r0_rd_out[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5237.490 0.000 5237.630 0.350 ;
    END
  END r0_rd_out[474]
  PIN r0_rd_out[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5248.530 0.000 5248.670 0.350 ;
    END
  END r0_rd_out[475]
  PIN r0_rd_out[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5259.570 0.000 5259.710 0.350 ;
    END
  END r0_rd_out[476]
  PIN r0_rd_out[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5270.610 0.000 5270.750 0.350 ;
    END
  END r0_rd_out[477]
  PIN r0_rd_out[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5281.650 0.000 5281.790 0.350 ;
    END
  END r0_rd_out[478]
  PIN r0_rd_out[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5292.690 0.000 5292.830 0.350 ;
    END
  END r0_rd_out[479]
  PIN r0_rd_out[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5303.730 0.000 5303.870 0.350 ;
    END
  END r0_rd_out[480]
  PIN r0_rd_out[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5314.770 0.000 5314.910 0.350 ;
    END
  END r0_rd_out[481]
  PIN r0_rd_out[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5325.810 0.000 5325.950 0.350 ;
    END
  END r0_rd_out[482]
  PIN r0_rd_out[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5336.850 0.000 5336.990 0.350 ;
    END
  END r0_rd_out[483]
  PIN r0_rd_out[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5347.890 0.000 5348.030 0.350 ;
    END
  END r0_rd_out[484]
  PIN r0_rd_out[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5358.930 0.000 5359.070 0.350 ;
    END
  END r0_rd_out[485]
  PIN r0_rd_out[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5369.970 0.000 5370.110 0.350 ;
    END
  END r0_rd_out[486]
  PIN r0_rd_out[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5381.010 0.000 5381.150 0.350 ;
    END
  END r0_rd_out[487]
  PIN r0_rd_out[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5392.050 0.000 5392.190 0.350 ;
    END
  END r0_rd_out[488]
  PIN r0_rd_out[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5403.090 0.000 5403.230 0.350 ;
    END
  END r0_rd_out[489]
  PIN r0_rd_out[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5414.130 0.000 5414.270 0.350 ;
    END
  END r0_rd_out[490]
  PIN r0_rd_out[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5425.170 0.000 5425.310 0.350 ;
    END
  END r0_rd_out[491]
  PIN r0_rd_out[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5436.210 0.000 5436.350 0.350 ;
    END
  END r0_rd_out[492]
  PIN r0_rd_out[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5447.250 0.000 5447.390 0.350 ;
    END
  END r0_rd_out[493]
  PIN r0_rd_out[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5458.290 0.000 5458.430 0.350 ;
    END
  END r0_rd_out[494]
  PIN r0_rd_out[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5469.330 0.000 5469.470 0.350 ;
    END
  END r0_rd_out[495]
  PIN r0_rd_out[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5480.370 0.000 5480.510 0.350 ;
    END
  END r0_rd_out[496]
  PIN r0_rd_out[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5491.410 0.000 5491.550 0.350 ;
    END
  END r0_rd_out[497]
  PIN r0_rd_out[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5502.450 0.000 5502.590 0.350 ;
    END
  END r0_rd_out[498]
  PIN r0_rd_out[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5513.490 0.000 5513.630 0.350 ;
    END
  END r0_rd_out[499]
  PIN r0_rd_out[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5524.530 0.000 5524.670 0.350 ;
    END
  END r0_rd_out[500]
  PIN r0_rd_out[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5535.570 0.000 5535.710 0.350 ;
    END
  END r0_rd_out[501]
  PIN r0_rd_out[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5546.610 0.000 5546.750 0.350 ;
    END
  END r0_rd_out[502]
  PIN r0_rd_out[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5557.650 0.000 5557.790 0.350 ;
    END
  END r0_rd_out[503]
  PIN r0_rd_out[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5568.690 0.000 5568.830 0.350 ;
    END
  END r0_rd_out[504]
  PIN r0_rd_out[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5579.730 0.000 5579.870 0.350 ;
    END
  END r0_rd_out[505]
  PIN r0_rd_out[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5590.770 0.000 5590.910 0.350 ;
    END
  END r0_rd_out[506]
  PIN r0_rd_out[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5601.810 0.000 5601.950 0.350 ;
    END
  END r0_rd_out[507]
  PIN r0_rd_out[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5612.850 0.000 5612.990 0.350 ;
    END
  END r0_rd_out[508]
  PIN r0_rd_out[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5623.890 0.000 5624.030 0.350 ;
    END
  END r0_rd_out[509]
  PIN r0_rd_out[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5634.930 0.000 5635.070 0.350 ;
    END
  END r0_rd_out[510]
  PIN r0_rd_out[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 5645.970 0.000 5646.110 0.350 ;
    END
  END r0_rd_out[511]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 6.650 5871.900 6.950 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 9.370 5871.900 9.670 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 12.090 5871.900 12.390 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 14.810 5871.900 15.110 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 17.530 5871.900 17.830 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 20.250 5871.900 20.550 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 22.970 5871.900 23.270 ;
    END
  END w0_addr_in[6]
  PIN w0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 25.690 5871.900 25.990 ;
    END
  END w0_addr_in[7]
  PIN w0_addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 28.410 5871.900 28.710 ;
    END
  END w0_addr_in[8]
  PIN w0_addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 31.130 5871.900 31.430 ;
    END
  END w0_addr_in[9]
  PIN w0_addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 33.850 5871.900 34.150 ;
    END
  END w0_addr_in[10]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 1435.810 4.670 1436.160 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 15.570 1435.810 15.710 1436.160 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 26.610 1435.810 26.750 1436.160 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 37.650 1435.810 37.790 1436.160 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 48.690 1435.810 48.830 1436.160 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 59.730 1435.810 59.870 1436.160 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 70.770 1435.810 70.910 1436.160 ;
    END
  END r0_addr_in[6]
  PIN r0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 81.810 1435.810 81.950 1436.160 ;
    END
  END r0_addr_in[7]
  PIN r0_addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 92.850 1435.810 92.990 1436.160 ;
    END
  END r0_addr_in[8]
  PIN r0_addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 103.890 1435.810 104.030 1436.160 ;
    END
  END r0_addr_in[9]
  PIN r0_addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 114.930 1435.810 115.070 1436.160 ;
    END
  END r0_addr_in[10]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 44.730 5871.900 45.030 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 55.610 5871.900 55.910 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 5871.100 66.490 5871.900 66.790 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 208.770 1435.810 208.910 1436.160 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 302.610 1435.810 302.750 1436.160 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 3.240 6.800 5.960 1429.360 ;
      RECT 14.120 6.800 16.840 1429.360 ;
      RECT 25.000 6.800 27.720 1429.360 ;
      RECT 35.880 6.800 38.600 1429.360 ;
      RECT 46.760 6.800 49.480 1429.360 ;
      RECT 57.640 6.800 60.360 1429.360 ;
      RECT 68.520 6.800 71.240 1429.360 ;
      RECT 79.400 6.800 82.120 1429.360 ;
      RECT 90.280 6.800 93.000 1429.360 ;
      RECT 101.160 6.800 103.880 1429.360 ;
      RECT 112.040 6.800 114.760 1429.360 ;
      RECT 122.920 6.800 125.640 1429.360 ;
      RECT 133.800 6.800 136.520 1429.360 ;
      RECT 144.680 6.800 147.400 1429.360 ;
      RECT 155.560 6.800 158.280 1429.360 ;
      RECT 166.440 6.800 169.160 1429.360 ;
      RECT 177.320 6.800 180.040 1429.360 ;
      RECT 188.200 6.800 190.920 1429.360 ;
      RECT 199.080 6.800 201.800 1429.360 ;
      RECT 209.960 6.800 212.680 1429.360 ;
      RECT 220.840 6.800 223.560 1429.360 ;
      RECT 231.720 6.800 234.440 1429.360 ;
      RECT 242.600 6.800 245.320 1429.360 ;
      RECT 253.480 6.800 256.200 1429.360 ;
      RECT 264.360 6.800 267.080 1429.360 ;
      RECT 275.240 6.800 277.960 1429.360 ;
      RECT 286.120 6.800 288.840 1429.360 ;
      RECT 297.000 6.800 299.720 1429.360 ;
      RECT 307.880 6.800 310.600 1429.360 ;
      RECT 318.760 6.800 321.480 1429.360 ;
      RECT 329.640 6.800 332.360 1429.360 ;
      RECT 340.520 6.800 343.240 1429.360 ;
      RECT 351.400 6.800 354.120 1429.360 ;
      RECT 362.280 6.800 365.000 1429.360 ;
      RECT 373.160 6.800 375.880 1429.360 ;
      RECT 384.040 6.800 386.760 1429.360 ;
      RECT 394.920 6.800 397.640 1429.360 ;
      RECT 405.800 6.800 408.520 1429.360 ;
      RECT 416.680 6.800 419.400 1429.360 ;
      RECT 427.560 6.800 430.280 1429.360 ;
      RECT 438.440 6.800 441.160 1429.360 ;
      RECT 449.320 6.800 452.040 1429.360 ;
      RECT 460.200 6.800 462.920 1429.360 ;
      RECT 471.080 6.800 473.800 1429.360 ;
      RECT 481.960 6.800 484.680 1429.360 ;
      RECT 492.840 6.800 495.560 1429.360 ;
      RECT 503.720 6.800 506.440 1429.360 ;
      RECT 514.600 6.800 517.320 1429.360 ;
      RECT 525.480 6.800 528.200 1429.360 ;
      RECT 536.360 6.800 539.080 1429.360 ;
      RECT 547.240 6.800 549.960 1429.360 ;
      RECT 558.120 6.800 560.840 1429.360 ;
      RECT 569.000 6.800 571.720 1429.360 ;
      RECT 579.880 6.800 582.600 1429.360 ;
      RECT 590.760 6.800 593.480 1429.360 ;
      RECT 601.640 6.800 604.360 1429.360 ;
      RECT 612.520 6.800 615.240 1429.360 ;
      RECT 623.400 6.800 626.120 1429.360 ;
      RECT 634.280 6.800 637.000 1429.360 ;
      RECT 645.160 6.800 647.880 1429.360 ;
      RECT 656.040 6.800 658.760 1429.360 ;
      RECT 666.920 6.800 669.640 1429.360 ;
      RECT 677.800 6.800 680.520 1429.360 ;
      RECT 688.680 6.800 691.400 1429.360 ;
      RECT 699.560 6.800 702.280 1429.360 ;
      RECT 710.440 6.800 713.160 1429.360 ;
      RECT 721.320 6.800 724.040 1429.360 ;
      RECT 732.200 6.800 734.920 1429.360 ;
      RECT 743.080 6.800 745.800 1429.360 ;
      RECT 753.960 6.800 756.680 1429.360 ;
      RECT 764.840 6.800 767.560 1429.360 ;
      RECT 775.720 6.800 778.440 1429.360 ;
      RECT 786.600 6.800 789.320 1429.360 ;
      RECT 797.480 6.800 800.200 1429.360 ;
      RECT 808.360 6.800 811.080 1429.360 ;
      RECT 819.240 6.800 821.960 1429.360 ;
      RECT 830.120 6.800 832.840 1429.360 ;
      RECT 841.000 6.800 843.720 1429.360 ;
      RECT 851.880 6.800 854.600 1429.360 ;
      RECT 862.760 6.800 865.480 1429.360 ;
      RECT 873.640 6.800 876.360 1429.360 ;
      RECT 884.520 6.800 887.240 1429.360 ;
      RECT 895.400 6.800 898.120 1429.360 ;
      RECT 906.280 6.800 909.000 1429.360 ;
      RECT 917.160 6.800 919.880 1429.360 ;
      RECT 928.040 6.800 930.760 1429.360 ;
      RECT 938.920 6.800 941.640 1429.360 ;
      RECT 949.800 6.800 952.520 1429.360 ;
      RECT 960.680 6.800 963.400 1429.360 ;
      RECT 971.560 6.800 974.280 1429.360 ;
      RECT 982.440 6.800 985.160 1429.360 ;
      RECT 993.320 6.800 996.040 1429.360 ;
      RECT 1004.200 6.800 1006.920 1429.360 ;
      RECT 1015.080 6.800 1017.800 1429.360 ;
      RECT 1025.960 6.800 1028.680 1429.360 ;
      RECT 1036.840 6.800 1039.560 1429.360 ;
      RECT 1047.720 6.800 1050.440 1429.360 ;
      RECT 1058.600 6.800 1061.320 1429.360 ;
      RECT 1069.480 6.800 1072.200 1429.360 ;
      RECT 1080.360 6.800 1083.080 1429.360 ;
      RECT 1091.240 6.800 1093.960 1429.360 ;
      RECT 1102.120 6.800 1104.840 1429.360 ;
      RECT 1113.000 6.800 1115.720 1429.360 ;
      RECT 1123.880 6.800 1126.600 1429.360 ;
      RECT 1134.760 6.800 1137.480 1429.360 ;
      RECT 1145.640 6.800 1148.360 1429.360 ;
      RECT 1156.520 6.800 1159.240 1429.360 ;
      RECT 1167.400 6.800 1170.120 1429.360 ;
      RECT 1178.280 6.800 1181.000 1429.360 ;
      RECT 1189.160 6.800 1191.880 1429.360 ;
      RECT 1200.040 6.800 1202.760 1429.360 ;
      RECT 1210.920 6.800 1213.640 1429.360 ;
      RECT 1221.800 6.800 1224.520 1429.360 ;
      RECT 1232.680 6.800 1235.400 1429.360 ;
      RECT 1243.560 6.800 1246.280 1429.360 ;
      RECT 1254.440 6.800 1257.160 1429.360 ;
      RECT 1265.320 6.800 1268.040 1429.360 ;
      RECT 1276.200 6.800 1278.920 1429.360 ;
      RECT 1287.080 6.800 1289.800 1429.360 ;
      RECT 1297.960 6.800 1300.680 1429.360 ;
      RECT 1308.840 6.800 1311.560 1429.360 ;
      RECT 1319.720 6.800 1322.440 1429.360 ;
      RECT 1330.600 6.800 1333.320 1429.360 ;
      RECT 1341.480 6.800 1344.200 1429.360 ;
      RECT 1352.360 6.800 1355.080 1429.360 ;
      RECT 1363.240 6.800 1365.960 1429.360 ;
      RECT 1374.120 6.800 1376.840 1429.360 ;
      RECT 1385.000 6.800 1387.720 1429.360 ;
      RECT 1395.880 6.800 1398.600 1429.360 ;
      RECT 1406.760 6.800 1409.480 1429.360 ;
      RECT 1417.640 6.800 1420.360 1429.360 ;
      RECT 1428.520 6.800 1431.240 1429.360 ;
      RECT 1439.400 6.800 1442.120 1429.360 ;
      RECT 1450.280 6.800 1453.000 1429.360 ;
      RECT 1461.160 6.800 1463.880 1429.360 ;
      RECT 1472.040 6.800 1474.760 1429.360 ;
      RECT 1482.920 6.800 1485.640 1429.360 ;
      RECT 1493.800 6.800 1496.520 1429.360 ;
      RECT 1504.680 6.800 1507.400 1429.360 ;
      RECT 1515.560 6.800 1518.280 1429.360 ;
      RECT 1526.440 6.800 1529.160 1429.360 ;
      RECT 1537.320 6.800 1540.040 1429.360 ;
      RECT 1548.200 6.800 1550.920 1429.360 ;
      RECT 1559.080 6.800 1561.800 1429.360 ;
      RECT 1569.960 6.800 1572.680 1429.360 ;
      RECT 1580.840 6.800 1583.560 1429.360 ;
      RECT 1591.720 6.800 1594.440 1429.360 ;
      RECT 1602.600 6.800 1605.320 1429.360 ;
      RECT 1613.480 6.800 1616.200 1429.360 ;
      RECT 1624.360 6.800 1627.080 1429.360 ;
      RECT 1635.240 6.800 1637.960 1429.360 ;
      RECT 1646.120 6.800 1648.840 1429.360 ;
      RECT 1657.000 6.800 1659.720 1429.360 ;
      RECT 1667.880 6.800 1670.600 1429.360 ;
      RECT 1678.760 6.800 1681.480 1429.360 ;
      RECT 1689.640 6.800 1692.360 1429.360 ;
      RECT 1700.520 6.800 1703.240 1429.360 ;
      RECT 1711.400 6.800 1714.120 1429.360 ;
      RECT 1722.280 6.800 1725.000 1429.360 ;
      RECT 1733.160 6.800 1735.880 1429.360 ;
      RECT 1744.040 6.800 1746.760 1429.360 ;
      RECT 1754.920 6.800 1757.640 1429.360 ;
      RECT 1765.800 6.800 1768.520 1429.360 ;
      RECT 1776.680 6.800 1779.400 1429.360 ;
      RECT 1787.560 6.800 1790.280 1429.360 ;
      RECT 1798.440 6.800 1801.160 1429.360 ;
      RECT 1809.320 6.800 1812.040 1429.360 ;
      RECT 1820.200 6.800 1822.920 1429.360 ;
      RECT 1831.080 6.800 1833.800 1429.360 ;
      RECT 1841.960 6.800 1844.680 1429.360 ;
      RECT 1852.840 6.800 1855.560 1429.360 ;
      RECT 1863.720 6.800 1866.440 1429.360 ;
      RECT 1874.600 6.800 1877.320 1429.360 ;
      RECT 1885.480 6.800 1888.200 1429.360 ;
      RECT 1896.360 6.800 1899.080 1429.360 ;
      RECT 1907.240 6.800 1909.960 1429.360 ;
      RECT 1918.120 6.800 1920.840 1429.360 ;
      RECT 1929.000 6.800 1931.720 1429.360 ;
      RECT 1939.880 6.800 1942.600 1429.360 ;
      RECT 1950.760 6.800 1953.480 1429.360 ;
      RECT 1961.640 6.800 1964.360 1429.360 ;
      RECT 1972.520 6.800 1975.240 1429.360 ;
      RECT 1983.400 6.800 1986.120 1429.360 ;
      RECT 1994.280 6.800 1997.000 1429.360 ;
      RECT 2005.160 6.800 2007.880 1429.360 ;
      RECT 2016.040 6.800 2018.760 1429.360 ;
      RECT 2026.920 6.800 2029.640 1429.360 ;
      RECT 2037.800 6.800 2040.520 1429.360 ;
      RECT 2048.680 6.800 2051.400 1429.360 ;
      RECT 2059.560 6.800 2062.280 1429.360 ;
      RECT 2070.440 6.800 2073.160 1429.360 ;
      RECT 2081.320 6.800 2084.040 1429.360 ;
      RECT 2092.200 6.800 2094.920 1429.360 ;
      RECT 2103.080 6.800 2105.800 1429.360 ;
      RECT 2113.960 6.800 2116.680 1429.360 ;
      RECT 2124.840 6.800 2127.560 1429.360 ;
      RECT 2135.720 6.800 2138.440 1429.360 ;
      RECT 2146.600 6.800 2149.320 1429.360 ;
      RECT 2157.480 6.800 2160.200 1429.360 ;
      RECT 2168.360 6.800 2171.080 1429.360 ;
      RECT 2179.240 6.800 2181.960 1429.360 ;
      RECT 2190.120 6.800 2192.840 1429.360 ;
      RECT 2201.000 6.800 2203.720 1429.360 ;
      RECT 2211.880 6.800 2214.600 1429.360 ;
      RECT 2222.760 6.800 2225.480 1429.360 ;
      RECT 2233.640 6.800 2236.360 1429.360 ;
      RECT 2244.520 6.800 2247.240 1429.360 ;
      RECT 2255.400 6.800 2258.120 1429.360 ;
      RECT 2266.280 6.800 2269.000 1429.360 ;
      RECT 2277.160 6.800 2279.880 1429.360 ;
      RECT 2288.040 6.800 2290.760 1429.360 ;
      RECT 2298.920 6.800 2301.640 1429.360 ;
      RECT 2309.800 6.800 2312.520 1429.360 ;
      RECT 2320.680 6.800 2323.400 1429.360 ;
      RECT 2331.560 6.800 2334.280 1429.360 ;
      RECT 2342.440 6.800 2345.160 1429.360 ;
      RECT 2353.320 6.800 2356.040 1429.360 ;
      RECT 2364.200 6.800 2366.920 1429.360 ;
      RECT 2375.080 6.800 2377.800 1429.360 ;
      RECT 2385.960 6.800 2388.680 1429.360 ;
      RECT 2396.840 6.800 2399.560 1429.360 ;
      RECT 2407.720 6.800 2410.440 1429.360 ;
      RECT 2418.600 6.800 2421.320 1429.360 ;
      RECT 2429.480 6.800 2432.200 1429.360 ;
      RECT 2440.360 6.800 2443.080 1429.360 ;
      RECT 2451.240 6.800 2453.960 1429.360 ;
      RECT 2462.120 6.800 2464.840 1429.360 ;
      RECT 2473.000 6.800 2475.720 1429.360 ;
      RECT 2483.880 6.800 2486.600 1429.360 ;
      RECT 2494.760 6.800 2497.480 1429.360 ;
      RECT 2505.640 6.800 2508.360 1429.360 ;
      RECT 2516.520 6.800 2519.240 1429.360 ;
      RECT 2527.400 6.800 2530.120 1429.360 ;
      RECT 2538.280 6.800 2541.000 1429.360 ;
      RECT 2549.160 6.800 2551.880 1429.360 ;
      RECT 2560.040 6.800 2562.760 1429.360 ;
      RECT 2570.920 6.800 2573.640 1429.360 ;
      RECT 2581.800 6.800 2584.520 1429.360 ;
      RECT 2592.680 6.800 2595.400 1429.360 ;
      RECT 2603.560 6.800 2606.280 1429.360 ;
      RECT 2614.440 6.800 2617.160 1429.360 ;
      RECT 2625.320 6.800 2628.040 1429.360 ;
      RECT 2636.200 6.800 2638.920 1429.360 ;
      RECT 2647.080 6.800 2649.800 1429.360 ;
      RECT 2657.960 6.800 2660.680 1429.360 ;
      RECT 2668.840 6.800 2671.560 1429.360 ;
      RECT 2679.720 6.800 2682.440 1429.360 ;
      RECT 2690.600 6.800 2693.320 1429.360 ;
      RECT 2701.480 6.800 2704.200 1429.360 ;
      RECT 2712.360 6.800 2715.080 1429.360 ;
      RECT 2723.240 6.800 2725.960 1429.360 ;
      RECT 2734.120 6.800 2736.840 1429.360 ;
      RECT 2745.000 6.800 2747.720 1429.360 ;
      RECT 2755.880 6.800 2758.600 1429.360 ;
      RECT 2766.760 6.800 2769.480 1429.360 ;
      RECT 2777.640 6.800 2780.360 1429.360 ;
      RECT 2788.520 6.800 2791.240 1429.360 ;
      RECT 2799.400 6.800 2802.120 1429.360 ;
      RECT 2810.280 6.800 2813.000 1429.360 ;
      RECT 2821.160 6.800 2823.880 1429.360 ;
      RECT 2832.040 6.800 2834.760 1429.360 ;
      RECT 2842.920 6.800 2845.640 1429.360 ;
      RECT 2853.800 6.800 2856.520 1429.360 ;
      RECT 2864.680 6.800 2867.400 1429.360 ;
      RECT 2875.560 6.800 2878.280 1429.360 ;
      RECT 2886.440 6.800 2889.160 1429.360 ;
      RECT 2897.320 6.800 2900.040 1429.360 ;
      RECT 2908.200 6.800 2910.920 1429.360 ;
      RECT 2919.080 6.800 2921.800 1429.360 ;
      RECT 2929.960 6.800 2932.680 1429.360 ;
      RECT 2940.840 6.800 2943.560 1429.360 ;
      RECT 2951.720 6.800 2954.440 1429.360 ;
      RECT 2962.600 6.800 2965.320 1429.360 ;
      RECT 2973.480 6.800 2976.200 1429.360 ;
      RECT 2984.360 6.800 2987.080 1429.360 ;
      RECT 2995.240 6.800 2997.960 1429.360 ;
      RECT 3006.120 6.800 3008.840 1429.360 ;
      RECT 3017.000 6.800 3019.720 1429.360 ;
      RECT 3027.880 6.800 3030.600 1429.360 ;
      RECT 3038.760 6.800 3041.480 1429.360 ;
      RECT 3049.640 6.800 3052.360 1429.360 ;
      RECT 3060.520 6.800 3063.240 1429.360 ;
      RECT 3071.400 6.800 3074.120 1429.360 ;
      RECT 3082.280 6.800 3085.000 1429.360 ;
      RECT 3093.160 6.800 3095.880 1429.360 ;
      RECT 3104.040 6.800 3106.760 1429.360 ;
      RECT 3114.920 6.800 3117.640 1429.360 ;
      RECT 3125.800 6.800 3128.520 1429.360 ;
      RECT 3136.680 6.800 3139.400 1429.360 ;
      RECT 3147.560 6.800 3150.280 1429.360 ;
      RECT 3158.440 6.800 3161.160 1429.360 ;
      RECT 3169.320 6.800 3172.040 1429.360 ;
      RECT 3180.200 6.800 3182.920 1429.360 ;
      RECT 3191.080 6.800 3193.800 1429.360 ;
      RECT 3201.960 6.800 3204.680 1429.360 ;
      RECT 3212.840 6.800 3215.560 1429.360 ;
      RECT 3223.720 6.800 3226.440 1429.360 ;
      RECT 3234.600 6.800 3237.320 1429.360 ;
      RECT 3245.480 6.800 3248.200 1429.360 ;
      RECT 3256.360 6.800 3259.080 1429.360 ;
      RECT 3267.240 6.800 3269.960 1429.360 ;
      RECT 3278.120 6.800 3280.840 1429.360 ;
      RECT 3289.000 6.800 3291.720 1429.360 ;
      RECT 3299.880 6.800 3302.600 1429.360 ;
      RECT 3310.760 6.800 3313.480 1429.360 ;
      RECT 3321.640 6.800 3324.360 1429.360 ;
      RECT 3332.520 6.800 3335.240 1429.360 ;
      RECT 3343.400 6.800 3346.120 1429.360 ;
      RECT 3354.280 6.800 3357.000 1429.360 ;
      RECT 3365.160 6.800 3367.880 1429.360 ;
      RECT 3376.040 6.800 3378.760 1429.360 ;
      RECT 3386.920 6.800 3389.640 1429.360 ;
      RECT 3397.800 6.800 3400.520 1429.360 ;
      RECT 3408.680 6.800 3411.400 1429.360 ;
      RECT 3419.560 6.800 3422.280 1429.360 ;
      RECT 3430.440 6.800 3433.160 1429.360 ;
      RECT 3441.320 6.800 3444.040 1429.360 ;
      RECT 3452.200 6.800 3454.920 1429.360 ;
      RECT 3463.080 6.800 3465.800 1429.360 ;
      RECT 3473.960 6.800 3476.680 1429.360 ;
      RECT 3484.840 6.800 3487.560 1429.360 ;
      RECT 3495.720 6.800 3498.440 1429.360 ;
      RECT 3506.600 6.800 3509.320 1429.360 ;
      RECT 3517.480 6.800 3520.200 1429.360 ;
      RECT 3528.360 6.800 3531.080 1429.360 ;
      RECT 3539.240 6.800 3541.960 1429.360 ;
      RECT 3550.120 6.800 3552.840 1429.360 ;
      RECT 3561.000 6.800 3563.720 1429.360 ;
      RECT 3571.880 6.800 3574.600 1429.360 ;
      RECT 3582.760 6.800 3585.480 1429.360 ;
      RECT 3593.640 6.800 3596.360 1429.360 ;
      RECT 3604.520 6.800 3607.240 1429.360 ;
      RECT 3615.400 6.800 3618.120 1429.360 ;
      RECT 3626.280 6.800 3629.000 1429.360 ;
      RECT 3637.160 6.800 3639.880 1429.360 ;
      RECT 3648.040 6.800 3650.760 1429.360 ;
      RECT 3658.920 6.800 3661.640 1429.360 ;
      RECT 3669.800 6.800 3672.520 1429.360 ;
      RECT 3680.680 6.800 3683.400 1429.360 ;
      RECT 3691.560 6.800 3694.280 1429.360 ;
      RECT 3702.440 6.800 3705.160 1429.360 ;
      RECT 3713.320 6.800 3716.040 1429.360 ;
      RECT 3724.200 6.800 3726.920 1429.360 ;
      RECT 3735.080 6.800 3737.800 1429.360 ;
      RECT 3745.960 6.800 3748.680 1429.360 ;
      RECT 3756.840 6.800 3759.560 1429.360 ;
      RECT 3767.720 6.800 3770.440 1429.360 ;
      RECT 3778.600 6.800 3781.320 1429.360 ;
      RECT 3789.480 6.800 3792.200 1429.360 ;
      RECT 3800.360 6.800 3803.080 1429.360 ;
      RECT 3811.240 6.800 3813.960 1429.360 ;
      RECT 3822.120 6.800 3824.840 1429.360 ;
      RECT 3833.000 6.800 3835.720 1429.360 ;
      RECT 3843.880 6.800 3846.600 1429.360 ;
      RECT 3854.760 6.800 3857.480 1429.360 ;
      RECT 3865.640 6.800 3868.360 1429.360 ;
      RECT 3876.520 6.800 3879.240 1429.360 ;
      RECT 3887.400 6.800 3890.120 1429.360 ;
      RECT 3898.280 6.800 3901.000 1429.360 ;
      RECT 3909.160 6.800 3911.880 1429.360 ;
      RECT 3920.040 6.800 3922.760 1429.360 ;
      RECT 3930.920 6.800 3933.640 1429.360 ;
      RECT 3941.800 6.800 3944.520 1429.360 ;
      RECT 3952.680 6.800 3955.400 1429.360 ;
      RECT 3963.560 6.800 3966.280 1429.360 ;
      RECT 3974.440 6.800 3977.160 1429.360 ;
      RECT 3985.320 6.800 3988.040 1429.360 ;
      RECT 3996.200 6.800 3998.920 1429.360 ;
      RECT 4007.080 6.800 4009.800 1429.360 ;
      RECT 4017.960 6.800 4020.680 1429.360 ;
      RECT 4028.840 6.800 4031.560 1429.360 ;
      RECT 4039.720 6.800 4042.440 1429.360 ;
      RECT 4050.600 6.800 4053.320 1429.360 ;
      RECT 4061.480 6.800 4064.200 1429.360 ;
      RECT 4072.360 6.800 4075.080 1429.360 ;
      RECT 4083.240 6.800 4085.960 1429.360 ;
      RECT 4094.120 6.800 4096.840 1429.360 ;
      RECT 4105.000 6.800 4107.720 1429.360 ;
      RECT 4115.880 6.800 4118.600 1429.360 ;
      RECT 4126.760 6.800 4129.480 1429.360 ;
      RECT 4137.640 6.800 4140.360 1429.360 ;
      RECT 4148.520 6.800 4151.240 1429.360 ;
      RECT 4159.400 6.800 4162.120 1429.360 ;
      RECT 4170.280 6.800 4173.000 1429.360 ;
      RECT 4181.160 6.800 4183.880 1429.360 ;
      RECT 4192.040 6.800 4194.760 1429.360 ;
      RECT 4202.920 6.800 4205.640 1429.360 ;
      RECT 4213.800 6.800 4216.520 1429.360 ;
      RECT 4224.680 6.800 4227.400 1429.360 ;
      RECT 4235.560 6.800 4238.280 1429.360 ;
      RECT 4246.440 6.800 4249.160 1429.360 ;
      RECT 4257.320 6.800 4260.040 1429.360 ;
      RECT 4268.200 6.800 4270.920 1429.360 ;
      RECT 4279.080 6.800 4281.800 1429.360 ;
      RECT 4289.960 6.800 4292.680 1429.360 ;
      RECT 4300.840 6.800 4303.560 1429.360 ;
      RECT 4311.720 6.800 4314.440 1429.360 ;
      RECT 4322.600 6.800 4325.320 1429.360 ;
      RECT 4333.480 6.800 4336.200 1429.360 ;
      RECT 4344.360 6.800 4347.080 1429.360 ;
      RECT 4355.240 6.800 4357.960 1429.360 ;
      RECT 4366.120 6.800 4368.840 1429.360 ;
      RECT 4377.000 6.800 4379.720 1429.360 ;
      RECT 4387.880 6.800 4390.600 1429.360 ;
      RECT 4398.760 6.800 4401.480 1429.360 ;
      RECT 4409.640 6.800 4412.360 1429.360 ;
      RECT 4420.520 6.800 4423.240 1429.360 ;
      RECT 4431.400 6.800 4434.120 1429.360 ;
      RECT 4442.280 6.800 4445.000 1429.360 ;
      RECT 4453.160 6.800 4455.880 1429.360 ;
      RECT 4464.040 6.800 4466.760 1429.360 ;
      RECT 4474.920 6.800 4477.640 1429.360 ;
      RECT 4485.800 6.800 4488.520 1429.360 ;
      RECT 4496.680 6.800 4499.400 1429.360 ;
      RECT 4507.560 6.800 4510.280 1429.360 ;
      RECT 4518.440 6.800 4521.160 1429.360 ;
      RECT 4529.320 6.800 4532.040 1429.360 ;
      RECT 4540.200 6.800 4542.920 1429.360 ;
      RECT 4551.080 6.800 4553.800 1429.360 ;
      RECT 4561.960 6.800 4564.680 1429.360 ;
      RECT 4572.840 6.800 4575.560 1429.360 ;
      RECT 4583.720 6.800 4586.440 1429.360 ;
      RECT 4594.600 6.800 4597.320 1429.360 ;
      RECT 4605.480 6.800 4608.200 1429.360 ;
      RECT 4616.360 6.800 4619.080 1429.360 ;
      RECT 4627.240 6.800 4629.960 1429.360 ;
      RECT 4638.120 6.800 4640.840 1429.360 ;
      RECT 4649.000 6.800 4651.720 1429.360 ;
      RECT 4659.880 6.800 4662.600 1429.360 ;
      RECT 4670.760 6.800 4673.480 1429.360 ;
      RECT 4681.640 6.800 4684.360 1429.360 ;
      RECT 4692.520 6.800 4695.240 1429.360 ;
      RECT 4703.400 6.800 4706.120 1429.360 ;
      RECT 4714.280 6.800 4717.000 1429.360 ;
      RECT 4725.160 6.800 4727.880 1429.360 ;
      RECT 4736.040 6.800 4738.760 1429.360 ;
      RECT 4746.920 6.800 4749.640 1429.360 ;
      RECT 4757.800 6.800 4760.520 1429.360 ;
      RECT 4768.680 6.800 4771.400 1429.360 ;
      RECT 4779.560 6.800 4782.280 1429.360 ;
      RECT 4790.440 6.800 4793.160 1429.360 ;
      RECT 4801.320 6.800 4804.040 1429.360 ;
      RECT 4812.200 6.800 4814.920 1429.360 ;
      RECT 4823.080 6.800 4825.800 1429.360 ;
      RECT 4833.960 6.800 4836.680 1429.360 ;
      RECT 4844.840 6.800 4847.560 1429.360 ;
      RECT 4855.720 6.800 4858.440 1429.360 ;
      RECT 4866.600 6.800 4869.320 1429.360 ;
      RECT 4877.480 6.800 4880.200 1429.360 ;
      RECT 4888.360 6.800 4891.080 1429.360 ;
      RECT 4899.240 6.800 4901.960 1429.360 ;
      RECT 4910.120 6.800 4912.840 1429.360 ;
      RECT 4921.000 6.800 4923.720 1429.360 ;
      RECT 4931.880 6.800 4934.600 1429.360 ;
      RECT 4942.760 6.800 4945.480 1429.360 ;
      RECT 4953.640 6.800 4956.360 1429.360 ;
      RECT 4964.520 6.800 4967.240 1429.360 ;
      RECT 4975.400 6.800 4978.120 1429.360 ;
      RECT 4986.280 6.800 4989.000 1429.360 ;
      RECT 4997.160 6.800 4999.880 1429.360 ;
      RECT 5008.040 6.800 5010.760 1429.360 ;
      RECT 5018.920 6.800 5021.640 1429.360 ;
      RECT 5029.800 6.800 5032.520 1429.360 ;
      RECT 5040.680 6.800 5043.400 1429.360 ;
      RECT 5051.560 6.800 5054.280 1429.360 ;
      RECT 5062.440 6.800 5065.160 1429.360 ;
      RECT 5073.320 6.800 5076.040 1429.360 ;
      RECT 5084.200 6.800 5086.920 1429.360 ;
      RECT 5095.080 6.800 5097.800 1429.360 ;
      RECT 5105.960 6.800 5108.680 1429.360 ;
      RECT 5116.840 6.800 5119.560 1429.360 ;
      RECT 5127.720 6.800 5130.440 1429.360 ;
      RECT 5138.600 6.800 5141.320 1429.360 ;
      RECT 5149.480 6.800 5152.200 1429.360 ;
      RECT 5160.360 6.800 5163.080 1429.360 ;
      RECT 5171.240 6.800 5173.960 1429.360 ;
      RECT 5182.120 6.800 5184.840 1429.360 ;
      RECT 5193.000 6.800 5195.720 1429.360 ;
      RECT 5203.880 6.800 5206.600 1429.360 ;
      RECT 5214.760 6.800 5217.480 1429.360 ;
      RECT 5225.640 6.800 5228.360 1429.360 ;
      RECT 5236.520 6.800 5239.240 1429.360 ;
      RECT 5247.400 6.800 5250.120 1429.360 ;
      RECT 5258.280 6.800 5261.000 1429.360 ;
      RECT 5269.160 6.800 5271.880 1429.360 ;
      RECT 5280.040 6.800 5282.760 1429.360 ;
      RECT 5290.920 6.800 5293.640 1429.360 ;
      RECT 5301.800 6.800 5304.520 1429.360 ;
      RECT 5312.680 6.800 5315.400 1429.360 ;
      RECT 5323.560 6.800 5326.280 1429.360 ;
      RECT 5334.440 6.800 5337.160 1429.360 ;
      RECT 5345.320 6.800 5348.040 1429.360 ;
      RECT 5356.200 6.800 5358.920 1429.360 ;
      RECT 5367.080 6.800 5369.800 1429.360 ;
      RECT 5377.960 6.800 5380.680 1429.360 ;
      RECT 5388.840 6.800 5391.560 1429.360 ;
      RECT 5399.720 6.800 5402.440 1429.360 ;
      RECT 5410.600 6.800 5413.320 1429.360 ;
      RECT 5421.480 6.800 5424.200 1429.360 ;
      RECT 5432.360 6.800 5435.080 1429.360 ;
      RECT 5443.240 6.800 5445.960 1429.360 ;
      RECT 5454.120 6.800 5456.840 1429.360 ;
      RECT 5465.000 6.800 5467.720 1429.360 ;
      RECT 5475.880 6.800 5478.600 1429.360 ;
      RECT 5486.760 6.800 5489.480 1429.360 ;
      RECT 5497.640 6.800 5500.360 1429.360 ;
      RECT 5508.520 6.800 5511.240 1429.360 ;
      RECT 5519.400 6.800 5522.120 1429.360 ;
      RECT 5530.280 6.800 5533.000 1429.360 ;
      RECT 5541.160 6.800 5543.880 1429.360 ;
      RECT 5552.040 6.800 5554.760 1429.360 ;
      RECT 5562.920 6.800 5565.640 1429.360 ;
      RECT 5573.800 6.800 5576.520 1429.360 ;
      RECT 5584.680 6.800 5587.400 1429.360 ;
      RECT 5595.560 6.800 5598.280 1429.360 ;
      RECT 5606.440 6.800 5609.160 1429.360 ;
      RECT 5617.320 6.800 5620.040 1429.360 ;
      RECT 5628.200 6.800 5630.920 1429.360 ;
      RECT 5639.080 6.800 5641.800 1429.360 ;
      RECT 5649.960 6.800 5652.680 1429.360 ;
      RECT 5660.840 6.800 5663.560 1429.360 ;
      RECT 5671.720 6.800 5674.440 1429.360 ;
      RECT 5682.600 6.800 5685.320 1429.360 ;
      RECT 5693.480 6.800 5696.200 1429.360 ;
      RECT 5704.360 6.800 5707.080 1429.360 ;
      RECT 5715.240 6.800 5717.960 1429.360 ;
      RECT 5726.120 6.800 5728.840 1429.360 ;
      RECT 5737.000 6.800 5739.720 1429.360 ;
      RECT 5747.880 6.800 5750.600 1429.360 ;
      RECT 5758.760 6.800 5761.480 1429.360 ;
      RECT 5769.640 6.800 5772.360 1429.360 ;
      RECT 5780.520 6.800 5783.240 1429.360 ;
      RECT 5791.400 6.800 5794.120 1429.360 ;
      RECT 5802.280 6.800 5805.000 1429.360 ;
      RECT 5813.160 6.800 5815.880 1429.360 ;
      RECT 5824.040 6.800 5826.760 1429.360 ;
      RECT 5834.920 6.800 5837.640 1429.360 ;
      RECT 5845.800 6.800 5848.520 1429.360 ;
      RECT 5856.680 6.800 5859.400 1429.360 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 8.680 6.800 11.400 1429.360 ;
      RECT 19.560 6.800 22.280 1429.360 ;
      RECT 30.440 6.800 33.160 1429.360 ;
      RECT 41.320 6.800 44.040 1429.360 ;
      RECT 52.200 6.800 54.920 1429.360 ;
      RECT 63.080 6.800 65.800 1429.360 ;
      RECT 73.960 6.800 76.680 1429.360 ;
      RECT 84.840 6.800 87.560 1429.360 ;
      RECT 95.720 6.800 98.440 1429.360 ;
      RECT 106.600 6.800 109.320 1429.360 ;
      RECT 117.480 6.800 120.200 1429.360 ;
      RECT 128.360 6.800 131.080 1429.360 ;
      RECT 139.240 6.800 141.960 1429.360 ;
      RECT 150.120 6.800 152.840 1429.360 ;
      RECT 161.000 6.800 163.720 1429.360 ;
      RECT 171.880 6.800 174.600 1429.360 ;
      RECT 182.760 6.800 185.480 1429.360 ;
      RECT 193.640 6.800 196.360 1429.360 ;
      RECT 204.520 6.800 207.240 1429.360 ;
      RECT 215.400 6.800 218.120 1429.360 ;
      RECT 226.280 6.800 229.000 1429.360 ;
      RECT 237.160 6.800 239.880 1429.360 ;
      RECT 248.040 6.800 250.760 1429.360 ;
      RECT 258.920 6.800 261.640 1429.360 ;
      RECT 269.800 6.800 272.520 1429.360 ;
      RECT 280.680 6.800 283.400 1429.360 ;
      RECT 291.560 6.800 294.280 1429.360 ;
      RECT 302.440 6.800 305.160 1429.360 ;
      RECT 313.320 6.800 316.040 1429.360 ;
      RECT 324.200 6.800 326.920 1429.360 ;
      RECT 335.080 6.800 337.800 1429.360 ;
      RECT 345.960 6.800 348.680 1429.360 ;
      RECT 356.840 6.800 359.560 1429.360 ;
      RECT 367.720 6.800 370.440 1429.360 ;
      RECT 378.600 6.800 381.320 1429.360 ;
      RECT 389.480 6.800 392.200 1429.360 ;
      RECT 400.360 6.800 403.080 1429.360 ;
      RECT 411.240 6.800 413.960 1429.360 ;
      RECT 422.120 6.800 424.840 1429.360 ;
      RECT 433.000 6.800 435.720 1429.360 ;
      RECT 443.880 6.800 446.600 1429.360 ;
      RECT 454.760 6.800 457.480 1429.360 ;
      RECT 465.640 6.800 468.360 1429.360 ;
      RECT 476.520 6.800 479.240 1429.360 ;
      RECT 487.400 6.800 490.120 1429.360 ;
      RECT 498.280 6.800 501.000 1429.360 ;
      RECT 509.160 6.800 511.880 1429.360 ;
      RECT 520.040 6.800 522.760 1429.360 ;
      RECT 530.920 6.800 533.640 1429.360 ;
      RECT 541.800 6.800 544.520 1429.360 ;
      RECT 552.680 6.800 555.400 1429.360 ;
      RECT 563.560 6.800 566.280 1429.360 ;
      RECT 574.440 6.800 577.160 1429.360 ;
      RECT 585.320 6.800 588.040 1429.360 ;
      RECT 596.200 6.800 598.920 1429.360 ;
      RECT 607.080 6.800 609.800 1429.360 ;
      RECT 617.960 6.800 620.680 1429.360 ;
      RECT 628.840 6.800 631.560 1429.360 ;
      RECT 639.720 6.800 642.440 1429.360 ;
      RECT 650.600 6.800 653.320 1429.360 ;
      RECT 661.480 6.800 664.200 1429.360 ;
      RECT 672.360 6.800 675.080 1429.360 ;
      RECT 683.240 6.800 685.960 1429.360 ;
      RECT 694.120 6.800 696.840 1429.360 ;
      RECT 705.000 6.800 707.720 1429.360 ;
      RECT 715.880 6.800 718.600 1429.360 ;
      RECT 726.760 6.800 729.480 1429.360 ;
      RECT 737.640 6.800 740.360 1429.360 ;
      RECT 748.520 6.800 751.240 1429.360 ;
      RECT 759.400 6.800 762.120 1429.360 ;
      RECT 770.280 6.800 773.000 1429.360 ;
      RECT 781.160 6.800 783.880 1429.360 ;
      RECT 792.040 6.800 794.760 1429.360 ;
      RECT 802.920 6.800 805.640 1429.360 ;
      RECT 813.800 6.800 816.520 1429.360 ;
      RECT 824.680 6.800 827.400 1429.360 ;
      RECT 835.560 6.800 838.280 1429.360 ;
      RECT 846.440 6.800 849.160 1429.360 ;
      RECT 857.320 6.800 860.040 1429.360 ;
      RECT 868.200 6.800 870.920 1429.360 ;
      RECT 879.080 6.800 881.800 1429.360 ;
      RECT 889.960 6.800 892.680 1429.360 ;
      RECT 900.840 6.800 903.560 1429.360 ;
      RECT 911.720 6.800 914.440 1429.360 ;
      RECT 922.600 6.800 925.320 1429.360 ;
      RECT 933.480 6.800 936.200 1429.360 ;
      RECT 944.360 6.800 947.080 1429.360 ;
      RECT 955.240 6.800 957.960 1429.360 ;
      RECT 966.120 6.800 968.840 1429.360 ;
      RECT 977.000 6.800 979.720 1429.360 ;
      RECT 987.880 6.800 990.600 1429.360 ;
      RECT 998.760 6.800 1001.480 1429.360 ;
      RECT 1009.640 6.800 1012.360 1429.360 ;
      RECT 1020.520 6.800 1023.240 1429.360 ;
      RECT 1031.400 6.800 1034.120 1429.360 ;
      RECT 1042.280 6.800 1045.000 1429.360 ;
      RECT 1053.160 6.800 1055.880 1429.360 ;
      RECT 1064.040 6.800 1066.760 1429.360 ;
      RECT 1074.920 6.800 1077.640 1429.360 ;
      RECT 1085.800 6.800 1088.520 1429.360 ;
      RECT 1096.680 6.800 1099.400 1429.360 ;
      RECT 1107.560 6.800 1110.280 1429.360 ;
      RECT 1118.440 6.800 1121.160 1429.360 ;
      RECT 1129.320 6.800 1132.040 1429.360 ;
      RECT 1140.200 6.800 1142.920 1429.360 ;
      RECT 1151.080 6.800 1153.800 1429.360 ;
      RECT 1161.960 6.800 1164.680 1429.360 ;
      RECT 1172.840 6.800 1175.560 1429.360 ;
      RECT 1183.720 6.800 1186.440 1429.360 ;
      RECT 1194.600 6.800 1197.320 1429.360 ;
      RECT 1205.480 6.800 1208.200 1429.360 ;
      RECT 1216.360 6.800 1219.080 1429.360 ;
      RECT 1227.240 6.800 1229.960 1429.360 ;
      RECT 1238.120 6.800 1240.840 1429.360 ;
      RECT 1249.000 6.800 1251.720 1429.360 ;
      RECT 1259.880 6.800 1262.600 1429.360 ;
      RECT 1270.760 6.800 1273.480 1429.360 ;
      RECT 1281.640 6.800 1284.360 1429.360 ;
      RECT 1292.520 6.800 1295.240 1429.360 ;
      RECT 1303.400 6.800 1306.120 1429.360 ;
      RECT 1314.280 6.800 1317.000 1429.360 ;
      RECT 1325.160 6.800 1327.880 1429.360 ;
      RECT 1336.040 6.800 1338.760 1429.360 ;
      RECT 1346.920 6.800 1349.640 1429.360 ;
      RECT 1357.800 6.800 1360.520 1429.360 ;
      RECT 1368.680 6.800 1371.400 1429.360 ;
      RECT 1379.560 6.800 1382.280 1429.360 ;
      RECT 1390.440 6.800 1393.160 1429.360 ;
      RECT 1401.320 6.800 1404.040 1429.360 ;
      RECT 1412.200 6.800 1414.920 1429.360 ;
      RECT 1423.080 6.800 1425.800 1429.360 ;
      RECT 1433.960 6.800 1436.680 1429.360 ;
      RECT 1444.840 6.800 1447.560 1429.360 ;
      RECT 1455.720 6.800 1458.440 1429.360 ;
      RECT 1466.600 6.800 1469.320 1429.360 ;
      RECT 1477.480 6.800 1480.200 1429.360 ;
      RECT 1488.360 6.800 1491.080 1429.360 ;
      RECT 1499.240 6.800 1501.960 1429.360 ;
      RECT 1510.120 6.800 1512.840 1429.360 ;
      RECT 1521.000 6.800 1523.720 1429.360 ;
      RECT 1531.880 6.800 1534.600 1429.360 ;
      RECT 1542.760 6.800 1545.480 1429.360 ;
      RECT 1553.640 6.800 1556.360 1429.360 ;
      RECT 1564.520 6.800 1567.240 1429.360 ;
      RECT 1575.400 6.800 1578.120 1429.360 ;
      RECT 1586.280 6.800 1589.000 1429.360 ;
      RECT 1597.160 6.800 1599.880 1429.360 ;
      RECT 1608.040 6.800 1610.760 1429.360 ;
      RECT 1618.920 6.800 1621.640 1429.360 ;
      RECT 1629.800 6.800 1632.520 1429.360 ;
      RECT 1640.680 6.800 1643.400 1429.360 ;
      RECT 1651.560 6.800 1654.280 1429.360 ;
      RECT 1662.440 6.800 1665.160 1429.360 ;
      RECT 1673.320 6.800 1676.040 1429.360 ;
      RECT 1684.200 6.800 1686.920 1429.360 ;
      RECT 1695.080 6.800 1697.800 1429.360 ;
      RECT 1705.960 6.800 1708.680 1429.360 ;
      RECT 1716.840 6.800 1719.560 1429.360 ;
      RECT 1727.720 6.800 1730.440 1429.360 ;
      RECT 1738.600 6.800 1741.320 1429.360 ;
      RECT 1749.480 6.800 1752.200 1429.360 ;
      RECT 1760.360 6.800 1763.080 1429.360 ;
      RECT 1771.240 6.800 1773.960 1429.360 ;
      RECT 1782.120 6.800 1784.840 1429.360 ;
      RECT 1793.000 6.800 1795.720 1429.360 ;
      RECT 1803.880 6.800 1806.600 1429.360 ;
      RECT 1814.760 6.800 1817.480 1429.360 ;
      RECT 1825.640 6.800 1828.360 1429.360 ;
      RECT 1836.520 6.800 1839.240 1429.360 ;
      RECT 1847.400 6.800 1850.120 1429.360 ;
      RECT 1858.280 6.800 1861.000 1429.360 ;
      RECT 1869.160 6.800 1871.880 1429.360 ;
      RECT 1880.040 6.800 1882.760 1429.360 ;
      RECT 1890.920 6.800 1893.640 1429.360 ;
      RECT 1901.800 6.800 1904.520 1429.360 ;
      RECT 1912.680 6.800 1915.400 1429.360 ;
      RECT 1923.560 6.800 1926.280 1429.360 ;
      RECT 1934.440 6.800 1937.160 1429.360 ;
      RECT 1945.320 6.800 1948.040 1429.360 ;
      RECT 1956.200 6.800 1958.920 1429.360 ;
      RECT 1967.080 6.800 1969.800 1429.360 ;
      RECT 1977.960 6.800 1980.680 1429.360 ;
      RECT 1988.840 6.800 1991.560 1429.360 ;
      RECT 1999.720 6.800 2002.440 1429.360 ;
      RECT 2010.600 6.800 2013.320 1429.360 ;
      RECT 2021.480 6.800 2024.200 1429.360 ;
      RECT 2032.360 6.800 2035.080 1429.360 ;
      RECT 2043.240 6.800 2045.960 1429.360 ;
      RECT 2054.120 6.800 2056.840 1429.360 ;
      RECT 2065.000 6.800 2067.720 1429.360 ;
      RECT 2075.880 6.800 2078.600 1429.360 ;
      RECT 2086.760 6.800 2089.480 1429.360 ;
      RECT 2097.640 6.800 2100.360 1429.360 ;
      RECT 2108.520 6.800 2111.240 1429.360 ;
      RECT 2119.400 6.800 2122.120 1429.360 ;
      RECT 2130.280 6.800 2133.000 1429.360 ;
      RECT 2141.160 6.800 2143.880 1429.360 ;
      RECT 2152.040 6.800 2154.760 1429.360 ;
      RECT 2162.920 6.800 2165.640 1429.360 ;
      RECT 2173.800 6.800 2176.520 1429.360 ;
      RECT 2184.680 6.800 2187.400 1429.360 ;
      RECT 2195.560 6.800 2198.280 1429.360 ;
      RECT 2206.440 6.800 2209.160 1429.360 ;
      RECT 2217.320 6.800 2220.040 1429.360 ;
      RECT 2228.200 6.800 2230.920 1429.360 ;
      RECT 2239.080 6.800 2241.800 1429.360 ;
      RECT 2249.960 6.800 2252.680 1429.360 ;
      RECT 2260.840 6.800 2263.560 1429.360 ;
      RECT 2271.720 6.800 2274.440 1429.360 ;
      RECT 2282.600 6.800 2285.320 1429.360 ;
      RECT 2293.480 6.800 2296.200 1429.360 ;
      RECT 2304.360 6.800 2307.080 1429.360 ;
      RECT 2315.240 6.800 2317.960 1429.360 ;
      RECT 2326.120 6.800 2328.840 1429.360 ;
      RECT 2337.000 6.800 2339.720 1429.360 ;
      RECT 2347.880 6.800 2350.600 1429.360 ;
      RECT 2358.760 6.800 2361.480 1429.360 ;
      RECT 2369.640 6.800 2372.360 1429.360 ;
      RECT 2380.520 6.800 2383.240 1429.360 ;
      RECT 2391.400 6.800 2394.120 1429.360 ;
      RECT 2402.280 6.800 2405.000 1429.360 ;
      RECT 2413.160 6.800 2415.880 1429.360 ;
      RECT 2424.040 6.800 2426.760 1429.360 ;
      RECT 2434.920 6.800 2437.640 1429.360 ;
      RECT 2445.800 6.800 2448.520 1429.360 ;
      RECT 2456.680 6.800 2459.400 1429.360 ;
      RECT 2467.560 6.800 2470.280 1429.360 ;
      RECT 2478.440 6.800 2481.160 1429.360 ;
      RECT 2489.320 6.800 2492.040 1429.360 ;
      RECT 2500.200 6.800 2502.920 1429.360 ;
      RECT 2511.080 6.800 2513.800 1429.360 ;
      RECT 2521.960 6.800 2524.680 1429.360 ;
      RECT 2532.840 6.800 2535.560 1429.360 ;
      RECT 2543.720 6.800 2546.440 1429.360 ;
      RECT 2554.600 6.800 2557.320 1429.360 ;
      RECT 2565.480 6.800 2568.200 1429.360 ;
      RECT 2576.360 6.800 2579.080 1429.360 ;
      RECT 2587.240 6.800 2589.960 1429.360 ;
      RECT 2598.120 6.800 2600.840 1429.360 ;
      RECT 2609.000 6.800 2611.720 1429.360 ;
      RECT 2619.880 6.800 2622.600 1429.360 ;
      RECT 2630.760 6.800 2633.480 1429.360 ;
      RECT 2641.640 6.800 2644.360 1429.360 ;
      RECT 2652.520 6.800 2655.240 1429.360 ;
      RECT 2663.400 6.800 2666.120 1429.360 ;
      RECT 2674.280 6.800 2677.000 1429.360 ;
      RECT 2685.160 6.800 2687.880 1429.360 ;
      RECT 2696.040 6.800 2698.760 1429.360 ;
      RECT 2706.920 6.800 2709.640 1429.360 ;
      RECT 2717.800 6.800 2720.520 1429.360 ;
      RECT 2728.680 6.800 2731.400 1429.360 ;
      RECT 2739.560 6.800 2742.280 1429.360 ;
      RECT 2750.440 6.800 2753.160 1429.360 ;
      RECT 2761.320 6.800 2764.040 1429.360 ;
      RECT 2772.200 6.800 2774.920 1429.360 ;
      RECT 2783.080 6.800 2785.800 1429.360 ;
      RECT 2793.960 6.800 2796.680 1429.360 ;
      RECT 2804.840 6.800 2807.560 1429.360 ;
      RECT 2815.720 6.800 2818.440 1429.360 ;
      RECT 2826.600 6.800 2829.320 1429.360 ;
      RECT 2837.480 6.800 2840.200 1429.360 ;
      RECT 2848.360 6.800 2851.080 1429.360 ;
      RECT 2859.240 6.800 2861.960 1429.360 ;
      RECT 2870.120 6.800 2872.840 1429.360 ;
      RECT 2881.000 6.800 2883.720 1429.360 ;
      RECT 2891.880 6.800 2894.600 1429.360 ;
      RECT 2902.760 6.800 2905.480 1429.360 ;
      RECT 2913.640 6.800 2916.360 1429.360 ;
      RECT 2924.520 6.800 2927.240 1429.360 ;
      RECT 2935.400 6.800 2938.120 1429.360 ;
      RECT 2946.280 6.800 2949.000 1429.360 ;
      RECT 2957.160 6.800 2959.880 1429.360 ;
      RECT 2968.040 6.800 2970.760 1429.360 ;
      RECT 2978.920 6.800 2981.640 1429.360 ;
      RECT 2989.800 6.800 2992.520 1429.360 ;
      RECT 3000.680 6.800 3003.400 1429.360 ;
      RECT 3011.560 6.800 3014.280 1429.360 ;
      RECT 3022.440 6.800 3025.160 1429.360 ;
      RECT 3033.320 6.800 3036.040 1429.360 ;
      RECT 3044.200 6.800 3046.920 1429.360 ;
      RECT 3055.080 6.800 3057.800 1429.360 ;
      RECT 3065.960 6.800 3068.680 1429.360 ;
      RECT 3076.840 6.800 3079.560 1429.360 ;
      RECT 3087.720 6.800 3090.440 1429.360 ;
      RECT 3098.600 6.800 3101.320 1429.360 ;
      RECT 3109.480 6.800 3112.200 1429.360 ;
      RECT 3120.360 6.800 3123.080 1429.360 ;
      RECT 3131.240 6.800 3133.960 1429.360 ;
      RECT 3142.120 6.800 3144.840 1429.360 ;
      RECT 3153.000 6.800 3155.720 1429.360 ;
      RECT 3163.880 6.800 3166.600 1429.360 ;
      RECT 3174.760 6.800 3177.480 1429.360 ;
      RECT 3185.640 6.800 3188.360 1429.360 ;
      RECT 3196.520 6.800 3199.240 1429.360 ;
      RECT 3207.400 6.800 3210.120 1429.360 ;
      RECT 3218.280 6.800 3221.000 1429.360 ;
      RECT 3229.160 6.800 3231.880 1429.360 ;
      RECT 3240.040 6.800 3242.760 1429.360 ;
      RECT 3250.920 6.800 3253.640 1429.360 ;
      RECT 3261.800 6.800 3264.520 1429.360 ;
      RECT 3272.680 6.800 3275.400 1429.360 ;
      RECT 3283.560 6.800 3286.280 1429.360 ;
      RECT 3294.440 6.800 3297.160 1429.360 ;
      RECT 3305.320 6.800 3308.040 1429.360 ;
      RECT 3316.200 6.800 3318.920 1429.360 ;
      RECT 3327.080 6.800 3329.800 1429.360 ;
      RECT 3337.960 6.800 3340.680 1429.360 ;
      RECT 3348.840 6.800 3351.560 1429.360 ;
      RECT 3359.720 6.800 3362.440 1429.360 ;
      RECT 3370.600 6.800 3373.320 1429.360 ;
      RECT 3381.480 6.800 3384.200 1429.360 ;
      RECT 3392.360 6.800 3395.080 1429.360 ;
      RECT 3403.240 6.800 3405.960 1429.360 ;
      RECT 3414.120 6.800 3416.840 1429.360 ;
      RECT 3425.000 6.800 3427.720 1429.360 ;
      RECT 3435.880 6.800 3438.600 1429.360 ;
      RECT 3446.760 6.800 3449.480 1429.360 ;
      RECT 3457.640 6.800 3460.360 1429.360 ;
      RECT 3468.520 6.800 3471.240 1429.360 ;
      RECT 3479.400 6.800 3482.120 1429.360 ;
      RECT 3490.280 6.800 3493.000 1429.360 ;
      RECT 3501.160 6.800 3503.880 1429.360 ;
      RECT 3512.040 6.800 3514.760 1429.360 ;
      RECT 3522.920 6.800 3525.640 1429.360 ;
      RECT 3533.800 6.800 3536.520 1429.360 ;
      RECT 3544.680 6.800 3547.400 1429.360 ;
      RECT 3555.560 6.800 3558.280 1429.360 ;
      RECT 3566.440 6.800 3569.160 1429.360 ;
      RECT 3577.320 6.800 3580.040 1429.360 ;
      RECT 3588.200 6.800 3590.920 1429.360 ;
      RECT 3599.080 6.800 3601.800 1429.360 ;
      RECT 3609.960 6.800 3612.680 1429.360 ;
      RECT 3620.840 6.800 3623.560 1429.360 ;
      RECT 3631.720 6.800 3634.440 1429.360 ;
      RECT 3642.600 6.800 3645.320 1429.360 ;
      RECT 3653.480 6.800 3656.200 1429.360 ;
      RECT 3664.360 6.800 3667.080 1429.360 ;
      RECT 3675.240 6.800 3677.960 1429.360 ;
      RECT 3686.120 6.800 3688.840 1429.360 ;
      RECT 3697.000 6.800 3699.720 1429.360 ;
      RECT 3707.880 6.800 3710.600 1429.360 ;
      RECT 3718.760 6.800 3721.480 1429.360 ;
      RECT 3729.640 6.800 3732.360 1429.360 ;
      RECT 3740.520 6.800 3743.240 1429.360 ;
      RECT 3751.400 6.800 3754.120 1429.360 ;
      RECT 3762.280 6.800 3765.000 1429.360 ;
      RECT 3773.160 6.800 3775.880 1429.360 ;
      RECT 3784.040 6.800 3786.760 1429.360 ;
      RECT 3794.920 6.800 3797.640 1429.360 ;
      RECT 3805.800 6.800 3808.520 1429.360 ;
      RECT 3816.680 6.800 3819.400 1429.360 ;
      RECT 3827.560 6.800 3830.280 1429.360 ;
      RECT 3838.440 6.800 3841.160 1429.360 ;
      RECT 3849.320 6.800 3852.040 1429.360 ;
      RECT 3860.200 6.800 3862.920 1429.360 ;
      RECT 3871.080 6.800 3873.800 1429.360 ;
      RECT 3881.960 6.800 3884.680 1429.360 ;
      RECT 3892.840 6.800 3895.560 1429.360 ;
      RECT 3903.720 6.800 3906.440 1429.360 ;
      RECT 3914.600 6.800 3917.320 1429.360 ;
      RECT 3925.480 6.800 3928.200 1429.360 ;
      RECT 3936.360 6.800 3939.080 1429.360 ;
      RECT 3947.240 6.800 3949.960 1429.360 ;
      RECT 3958.120 6.800 3960.840 1429.360 ;
      RECT 3969.000 6.800 3971.720 1429.360 ;
      RECT 3979.880 6.800 3982.600 1429.360 ;
      RECT 3990.760 6.800 3993.480 1429.360 ;
      RECT 4001.640 6.800 4004.360 1429.360 ;
      RECT 4012.520 6.800 4015.240 1429.360 ;
      RECT 4023.400 6.800 4026.120 1429.360 ;
      RECT 4034.280 6.800 4037.000 1429.360 ;
      RECT 4045.160 6.800 4047.880 1429.360 ;
      RECT 4056.040 6.800 4058.760 1429.360 ;
      RECT 4066.920 6.800 4069.640 1429.360 ;
      RECT 4077.800 6.800 4080.520 1429.360 ;
      RECT 4088.680 6.800 4091.400 1429.360 ;
      RECT 4099.560 6.800 4102.280 1429.360 ;
      RECT 4110.440 6.800 4113.160 1429.360 ;
      RECT 4121.320 6.800 4124.040 1429.360 ;
      RECT 4132.200 6.800 4134.920 1429.360 ;
      RECT 4143.080 6.800 4145.800 1429.360 ;
      RECT 4153.960 6.800 4156.680 1429.360 ;
      RECT 4164.840 6.800 4167.560 1429.360 ;
      RECT 4175.720 6.800 4178.440 1429.360 ;
      RECT 4186.600 6.800 4189.320 1429.360 ;
      RECT 4197.480 6.800 4200.200 1429.360 ;
      RECT 4208.360 6.800 4211.080 1429.360 ;
      RECT 4219.240 6.800 4221.960 1429.360 ;
      RECT 4230.120 6.800 4232.840 1429.360 ;
      RECT 4241.000 6.800 4243.720 1429.360 ;
      RECT 4251.880 6.800 4254.600 1429.360 ;
      RECT 4262.760 6.800 4265.480 1429.360 ;
      RECT 4273.640 6.800 4276.360 1429.360 ;
      RECT 4284.520 6.800 4287.240 1429.360 ;
      RECT 4295.400 6.800 4298.120 1429.360 ;
      RECT 4306.280 6.800 4309.000 1429.360 ;
      RECT 4317.160 6.800 4319.880 1429.360 ;
      RECT 4328.040 6.800 4330.760 1429.360 ;
      RECT 4338.920 6.800 4341.640 1429.360 ;
      RECT 4349.800 6.800 4352.520 1429.360 ;
      RECT 4360.680 6.800 4363.400 1429.360 ;
      RECT 4371.560 6.800 4374.280 1429.360 ;
      RECT 4382.440 6.800 4385.160 1429.360 ;
      RECT 4393.320 6.800 4396.040 1429.360 ;
      RECT 4404.200 6.800 4406.920 1429.360 ;
      RECT 4415.080 6.800 4417.800 1429.360 ;
      RECT 4425.960 6.800 4428.680 1429.360 ;
      RECT 4436.840 6.800 4439.560 1429.360 ;
      RECT 4447.720 6.800 4450.440 1429.360 ;
      RECT 4458.600 6.800 4461.320 1429.360 ;
      RECT 4469.480 6.800 4472.200 1429.360 ;
      RECT 4480.360 6.800 4483.080 1429.360 ;
      RECT 4491.240 6.800 4493.960 1429.360 ;
      RECT 4502.120 6.800 4504.840 1429.360 ;
      RECT 4513.000 6.800 4515.720 1429.360 ;
      RECT 4523.880 6.800 4526.600 1429.360 ;
      RECT 4534.760 6.800 4537.480 1429.360 ;
      RECT 4545.640 6.800 4548.360 1429.360 ;
      RECT 4556.520 6.800 4559.240 1429.360 ;
      RECT 4567.400 6.800 4570.120 1429.360 ;
      RECT 4578.280 6.800 4581.000 1429.360 ;
      RECT 4589.160 6.800 4591.880 1429.360 ;
      RECT 4600.040 6.800 4602.760 1429.360 ;
      RECT 4610.920 6.800 4613.640 1429.360 ;
      RECT 4621.800 6.800 4624.520 1429.360 ;
      RECT 4632.680 6.800 4635.400 1429.360 ;
      RECT 4643.560 6.800 4646.280 1429.360 ;
      RECT 4654.440 6.800 4657.160 1429.360 ;
      RECT 4665.320 6.800 4668.040 1429.360 ;
      RECT 4676.200 6.800 4678.920 1429.360 ;
      RECT 4687.080 6.800 4689.800 1429.360 ;
      RECT 4697.960 6.800 4700.680 1429.360 ;
      RECT 4708.840 6.800 4711.560 1429.360 ;
      RECT 4719.720 6.800 4722.440 1429.360 ;
      RECT 4730.600 6.800 4733.320 1429.360 ;
      RECT 4741.480 6.800 4744.200 1429.360 ;
      RECT 4752.360 6.800 4755.080 1429.360 ;
      RECT 4763.240 6.800 4765.960 1429.360 ;
      RECT 4774.120 6.800 4776.840 1429.360 ;
      RECT 4785.000 6.800 4787.720 1429.360 ;
      RECT 4795.880 6.800 4798.600 1429.360 ;
      RECT 4806.760 6.800 4809.480 1429.360 ;
      RECT 4817.640 6.800 4820.360 1429.360 ;
      RECT 4828.520 6.800 4831.240 1429.360 ;
      RECT 4839.400 6.800 4842.120 1429.360 ;
      RECT 4850.280 6.800 4853.000 1429.360 ;
      RECT 4861.160 6.800 4863.880 1429.360 ;
      RECT 4872.040 6.800 4874.760 1429.360 ;
      RECT 4882.920 6.800 4885.640 1429.360 ;
      RECT 4893.800 6.800 4896.520 1429.360 ;
      RECT 4904.680 6.800 4907.400 1429.360 ;
      RECT 4915.560 6.800 4918.280 1429.360 ;
      RECT 4926.440 6.800 4929.160 1429.360 ;
      RECT 4937.320 6.800 4940.040 1429.360 ;
      RECT 4948.200 6.800 4950.920 1429.360 ;
      RECT 4959.080 6.800 4961.800 1429.360 ;
      RECT 4969.960 6.800 4972.680 1429.360 ;
      RECT 4980.840 6.800 4983.560 1429.360 ;
      RECT 4991.720 6.800 4994.440 1429.360 ;
      RECT 5002.600 6.800 5005.320 1429.360 ;
      RECT 5013.480 6.800 5016.200 1429.360 ;
      RECT 5024.360 6.800 5027.080 1429.360 ;
      RECT 5035.240 6.800 5037.960 1429.360 ;
      RECT 5046.120 6.800 5048.840 1429.360 ;
      RECT 5057.000 6.800 5059.720 1429.360 ;
      RECT 5067.880 6.800 5070.600 1429.360 ;
      RECT 5078.760 6.800 5081.480 1429.360 ;
      RECT 5089.640 6.800 5092.360 1429.360 ;
      RECT 5100.520 6.800 5103.240 1429.360 ;
      RECT 5111.400 6.800 5114.120 1429.360 ;
      RECT 5122.280 6.800 5125.000 1429.360 ;
      RECT 5133.160 6.800 5135.880 1429.360 ;
      RECT 5144.040 6.800 5146.760 1429.360 ;
      RECT 5154.920 6.800 5157.640 1429.360 ;
      RECT 5165.800 6.800 5168.520 1429.360 ;
      RECT 5176.680 6.800 5179.400 1429.360 ;
      RECT 5187.560 6.800 5190.280 1429.360 ;
      RECT 5198.440 6.800 5201.160 1429.360 ;
      RECT 5209.320 6.800 5212.040 1429.360 ;
      RECT 5220.200 6.800 5222.920 1429.360 ;
      RECT 5231.080 6.800 5233.800 1429.360 ;
      RECT 5241.960 6.800 5244.680 1429.360 ;
      RECT 5252.840 6.800 5255.560 1429.360 ;
      RECT 5263.720 6.800 5266.440 1429.360 ;
      RECT 5274.600 6.800 5277.320 1429.360 ;
      RECT 5285.480 6.800 5288.200 1429.360 ;
      RECT 5296.360 6.800 5299.080 1429.360 ;
      RECT 5307.240 6.800 5309.960 1429.360 ;
      RECT 5318.120 6.800 5320.840 1429.360 ;
      RECT 5329.000 6.800 5331.720 1429.360 ;
      RECT 5339.880 6.800 5342.600 1429.360 ;
      RECT 5350.760 6.800 5353.480 1429.360 ;
      RECT 5361.640 6.800 5364.360 1429.360 ;
      RECT 5372.520 6.800 5375.240 1429.360 ;
      RECT 5383.400 6.800 5386.120 1429.360 ;
      RECT 5394.280 6.800 5397.000 1429.360 ;
      RECT 5405.160 6.800 5407.880 1429.360 ;
      RECT 5416.040 6.800 5418.760 1429.360 ;
      RECT 5426.920 6.800 5429.640 1429.360 ;
      RECT 5437.800 6.800 5440.520 1429.360 ;
      RECT 5448.680 6.800 5451.400 1429.360 ;
      RECT 5459.560 6.800 5462.280 1429.360 ;
      RECT 5470.440 6.800 5473.160 1429.360 ;
      RECT 5481.320 6.800 5484.040 1429.360 ;
      RECT 5492.200 6.800 5494.920 1429.360 ;
      RECT 5503.080 6.800 5505.800 1429.360 ;
      RECT 5513.960 6.800 5516.680 1429.360 ;
      RECT 5524.840 6.800 5527.560 1429.360 ;
      RECT 5535.720 6.800 5538.440 1429.360 ;
      RECT 5546.600 6.800 5549.320 1429.360 ;
      RECT 5557.480 6.800 5560.200 1429.360 ;
      RECT 5568.360 6.800 5571.080 1429.360 ;
      RECT 5579.240 6.800 5581.960 1429.360 ;
      RECT 5590.120 6.800 5592.840 1429.360 ;
      RECT 5601.000 6.800 5603.720 1429.360 ;
      RECT 5611.880 6.800 5614.600 1429.360 ;
      RECT 5622.760 6.800 5625.480 1429.360 ;
      RECT 5633.640 6.800 5636.360 1429.360 ;
      RECT 5644.520 6.800 5647.240 1429.360 ;
      RECT 5655.400 6.800 5658.120 1429.360 ;
      RECT 5666.280 6.800 5669.000 1429.360 ;
      RECT 5677.160 6.800 5679.880 1429.360 ;
      RECT 5688.040 6.800 5690.760 1429.360 ;
      RECT 5698.920 6.800 5701.640 1429.360 ;
      RECT 5709.800 6.800 5712.520 1429.360 ;
      RECT 5720.680 6.800 5723.400 1429.360 ;
      RECT 5731.560 6.800 5734.280 1429.360 ;
      RECT 5742.440 6.800 5745.160 1429.360 ;
      RECT 5753.320 6.800 5756.040 1429.360 ;
      RECT 5764.200 6.800 5766.920 1429.360 ;
      RECT 5775.080 6.800 5777.800 1429.360 ;
      RECT 5785.960 6.800 5788.680 1429.360 ;
      RECT 5796.840 6.800 5799.560 1429.360 ;
      RECT 5807.720 6.800 5810.440 1429.360 ;
      RECT 5818.600 6.800 5821.320 1429.360 ;
      RECT 5829.480 6.800 5832.200 1429.360 ;
      RECT 5840.360 6.800 5843.080 1429.360 ;
      RECT 5851.240 6.800 5853.960 1429.360 ;
      RECT 5862.120 6.800 5864.840 1429.360 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 5871.900 1436.160 ;
    LAYER met2 ;
    RECT 0 0 5871.900 1436.160 ;
    LAYER met3 ;
    RECT 0.800 0 5871.900 1436.160 ;
    LAYER met4 ;
    RECT 0 0 5871.900 6.800 ;
    RECT 0 1429.360 5871.900 1436.160 ;
    RECT 0.000 6.800 3.240 1429.360 ;
    RECT 5.960 6.800 8.680 1429.360 ;
    RECT 11.400 6.800 14.120 1429.360 ;
    RECT 16.840 6.800 19.560 1429.360 ;
    RECT 22.280 6.800 25.000 1429.360 ;
    RECT 27.720 6.800 30.440 1429.360 ;
    RECT 33.160 6.800 35.880 1429.360 ;
    RECT 38.600 6.800 41.320 1429.360 ;
    RECT 44.040 6.800 46.760 1429.360 ;
    RECT 49.480 6.800 52.200 1429.360 ;
    RECT 54.920 6.800 57.640 1429.360 ;
    RECT 60.360 6.800 63.080 1429.360 ;
    RECT 65.800 6.800 68.520 1429.360 ;
    RECT 71.240 6.800 73.960 1429.360 ;
    RECT 76.680 6.800 79.400 1429.360 ;
    RECT 82.120 6.800 84.840 1429.360 ;
    RECT 87.560 6.800 90.280 1429.360 ;
    RECT 93.000 6.800 95.720 1429.360 ;
    RECT 98.440 6.800 101.160 1429.360 ;
    RECT 103.880 6.800 106.600 1429.360 ;
    RECT 109.320 6.800 112.040 1429.360 ;
    RECT 114.760 6.800 117.480 1429.360 ;
    RECT 120.200 6.800 122.920 1429.360 ;
    RECT 125.640 6.800 128.360 1429.360 ;
    RECT 131.080 6.800 133.800 1429.360 ;
    RECT 136.520 6.800 139.240 1429.360 ;
    RECT 141.960 6.800 144.680 1429.360 ;
    RECT 147.400 6.800 150.120 1429.360 ;
    RECT 152.840 6.800 155.560 1429.360 ;
    RECT 158.280 6.800 161.000 1429.360 ;
    RECT 163.720 6.800 166.440 1429.360 ;
    RECT 169.160 6.800 171.880 1429.360 ;
    RECT 174.600 6.800 177.320 1429.360 ;
    RECT 180.040 6.800 182.760 1429.360 ;
    RECT 185.480 6.800 188.200 1429.360 ;
    RECT 190.920 6.800 193.640 1429.360 ;
    RECT 196.360 6.800 199.080 1429.360 ;
    RECT 201.800 6.800 204.520 1429.360 ;
    RECT 207.240 6.800 209.960 1429.360 ;
    RECT 212.680 6.800 215.400 1429.360 ;
    RECT 218.120 6.800 220.840 1429.360 ;
    RECT 223.560 6.800 226.280 1429.360 ;
    RECT 229.000 6.800 231.720 1429.360 ;
    RECT 234.440 6.800 237.160 1429.360 ;
    RECT 239.880 6.800 242.600 1429.360 ;
    RECT 245.320 6.800 248.040 1429.360 ;
    RECT 250.760 6.800 253.480 1429.360 ;
    RECT 256.200 6.800 258.920 1429.360 ;
    RECT 261.640 6.800 264.360 1429.360 ;
    RECT 267.080 6.800 269.800 1429.360 ;
    RECT 272.520 6.800 275.240 1429.360 ;
    RECT 277.960 6.800 280.680 1429.360 ;
    RECT 283.400 6.800 286.120 1429.360 ;
    RECT 288.840 6.800 291.560 1429.360 ;
    RECT 294.280 6.800 297.000 1429.360 ;
    RECT 299.720 6.800 302.440 1429.360 ;
    RECT 305.160 6.800 307.880 1429.360 ;
    RECT 310.600 6.800 313.320 1429.360 ;
    RECT 316.040 6.800 318.760 1429.360 ;
    RECT 321.480 6.800 324.200 1429.360 ;
    RECT 326.920 6.800 329.640 1429.360 ;
    RECT 332.360 6.800 335.080 1429.360 ;
    RECT 337.800 6.800 340.520 1429.360 ;
    RECT 343.240 6.800 345.960 1429.360 ;
    RECT 348.680 6.800 351.400 1429.360 ;
    RECT 354.120 6.800 356.840 1429.360 ;
    RECT 359.560 6.800 362.280 1429.360 ;
    RECT 365.000 6.800 367.720 1429.360 ;
    RECT 370.440 6.800 373.160 1429.360 ;
    RECT 375.880 6.800 378.600 1429.360 ;
    RECT 381.320 6.800 384.040 1429.360 ;
    RECT 386.760 6.800 389.480 1429.360 ;
    RECT 392.200 6.800 394.920 1429.360 ;
    RECT 397.640 6.800 400.360 1429.360 ;
    RECT 403.080 6.800 405.800 1429.360 ;
    RECT 408.520 6.800 411.240 1429.360 ;
    RECT 413.960 6.800 416.680 1429.360 ;
    RECT 419.400 6.800 422.120 1429.360 ;
    RECT 424.840 6.800 427.560 1429.360 ;
    RECT 430.280 6.800 433.000 1429.360 ;
    RECT 435.720 6.800 438.440 1429.360 ;
    RECT 441.160 6.800 443.880 1429.360 ;
    RECT 446.600 6.800 449.320 1429.360 ;
    RECT 452.040 6.800 454.760 1429.360 ;
    RECT 457.480 6.800 460.200 1429.360 ;
    RECT 462.920 6.800 465.640 1429.360 ;
    RECT 468.360 6.800 471.080 1429.360 ;
    RECT 473.800 6.800 476.520 1429.360 ;
    RECT 479.240 6.800 481.960 1429.360 ;
    RECT 484.680 6.800 487.400 1429.360 ;
    RECT 490.120 6.800 492.840 1429.360 ;
    RECT 495.560 6.800 498.280 1429.360 ;
    RECT 501.000 6.800 503.720 1429.360 ;
    RECT 506.440 6.800 509.160 1429.360 ;
    RECT 511.880 6.800 514.600 1429.360 ;
    RECT 517.320 6.800 520.040 1429.360 ;
    RECT 522.760 6.800 525.480 1429.360 ;
    RECT 528.200 6.800 530.920 1429.360 ;
    RECT 533.640 6.800 536.360 1429.360 ;
    RECT 539.080 6.800 541.800 1429.360 ;
    RECT 544.520 6.800 547.240 1429.360 ;
    RECT 549.960 6.800 552.680 1429.360 ;
    RECT 555.400 6.800 558.120 1429.360 ;
    RECT 560.840 6.800 563.560 1429.360 ;
    RECT 566.280 6.800 569.000 1429.360 ;
    RECT 571.720 6.800 574.440 1429.360 ;
    RECT 577.160 6.800 579.880 1429.360 ;
    RECT 582.600 6.800 585.320 1429.360 ;
    RECT 588.040 6.800 590.760 1429.360 ;
    RECT 593.480 6.800 596.200 1429.360 ;
    RECT 598.920 6.800 601.640 1429.360 ;
    RECT 604.360 6.800 607.080 1429.360 ;
    RECT 609.800 6.800 612.520 1429.360 ;
    RECT 615.240 6.800 617.960 1429.360 ;
    RECT 620.680 6.800 623.400 1429.360 ;
    RECT 626.120 6.800 628.840 1429.360 ;
    RECT 631.560 6.800 634.280 1429.360 ;
    RECT 637.000 6.800 639.720 1429.360 ;
    RECT 642.440 6.800 645.160 1429.360 ;
    RECT 647.880 6.800 650.600 1429.360 ;
    RECT 653.320 6.800 656.040 1429.360 ;
    RECT 658.760 6.800 661.480 1429.360 ;
    RECT 664.200 6.800 666.920 1429.360 ;
    RECT 669.640 6.800 672.360 1429.360 ;
    RECT 675.080 6.800 677.800 1429.360 ;
    RECT 680.520 6.800 683.240 1429.360 ;
    RECT 685.960 6.800 688.680 1429.360 ;
    RECT 691.400 6.800 694.120 1429.360 ;
    RECT 696.840 6.800 699.560 1429.360 ;
    RECT 702.280 6.800 705.000 1429.360 ;
    RECT 707.720 6.800 710.440 1429.360 ;
    RECT 713.160 6.800 715.880 1429.360 ;
    RECT 718.600 6.800 721.320 1429.360 ;
    RECT 724.040 6.800 726.760 1429.360 ;
    RECT 729.480 6.800 732.200 1429.360 ;
    RECT 734.920 6.800 737.640 1429.360 ;
    RECT 740.360 6.800 743.080 1429.360 ;
    RECT 745.800 6.800 748.520 1429.360 ;
    RECT 751.240 6.800 753.960 1429.360 ;
    RECT 756.680 6.800 759.400 1429.360 ;
    RECT 762.120 6.800 764.840 1429.360 ;
    RECT 767.560 6.800 770.280 1429.360 ;
    RECT 773.000 6.800 775.720 1429.360 ;
    RECT 778.440 6.800 781.160 1429.360 ;
    RECT 783.880 6.800 786.600 1429.360 ;
    RECT 789.320 6.800 792.040 1429.360 ;
    RECT 794.760 6.800 797.480 1429.360 ;
    RECT 800.200 6.800 802.920 1429.360 ;
    RECT 805.640 6.800 808.360 1429.360 ;
    RECT 811.080 6.800 813.800 1429.360 ;
    RECT 816.520 6.800 819.240 1429.360 ;
    RECT 821.960 6.800 824.680 1429.360 ;
    RECT 827.400 6.800 830.120 1429.360 ;
    RECT 832.840 6.800 835.560 1429.360 ;
    RECT 838.280 6.800 841.000 1429.360 ;
    RECT 843.720 6.800 846.440 1429.360 ;
    RECT 849.160 6.800 851.880 1429.360 ;
    RECT 854.600 6.800 857.320 1429.360 ;
    RECT 860.040 6.800 862.760 1429.360 ;
    RECT 865.480 6.800 868.200 1429.360 ;
    RECT 870.920 6.800 873.640 1429.360 ;
    RECT 876.360 6.800 879.080 1429.360 ;
    RECT 881.800 6.800 884.520 1429.360 ;
    RECT 887.240 6.800 889.960 1429.360 ;
    RECT 892.680 6.800 895.400 1429.360 ;
    RECT 898.120 6.800 900.840 1429.360 ;
    RECT 903.560 6.800 906.280 1429.360 ;
    RECT 909.000 6.800 911.720 1429.360 ;
    RECT 914.440 6.800 917.160 1429.360 ;
    RECT 919.880 6.800 922.600 1429.360 ;
    RECT 925.320 6.800 928.040 1429.360 ;
    RECT 930.760 6.800 933.480 1429.360 ;
    RECT 936.200 6.800 938.920 1429.360 ;
    RECT 941.640 6.800 944.360 1429.360 ;
    RECT 947.080 6.800 949.800 1429.360 ;
    RECT 952.520 6.800 955.240 1429.360 ;
    RECT 957.960 6.800 960.680 1429.360 ;
    RECT 963.400 6.800 966.120 1429.360 ;
    RECT 968.840 6.800 971.560 1429.360 ;
    RECT 974.280 6.800 977.000 1429.360 ;
    RECT 979.720 6.800 982.440 1429.360 ;
    RECT 985.160 6.800 987.880 1429.360 ;
    RECT 990.600 6.800 993.320 1429.360 ;
    RECT 996.040 6.800 998.760 1429.360 ;
    RECT 1001.480 6.800 1004.200 1429.360 ;
    RECT 1006.920 6.800 1009.640 1429.360 ;
    RECT 1012.360 6.800 1015.080 1429.360 ;
    RECT 1017.800 6.800 1020.520 1429.360 ;
    RECT 1023.240 6.800 1025.960 1429.360 ;
    RECT 1028.680 6.800 1031.400 1429.360 ;
    RECT 1034.120 6.800 1036.840 1429.360 ;
    RECT 1039.560 6.800 1042.280 1429.360 ;
    RECT 1045.000 6.800 1047.720 1429.360 ;
    RECT 1050.440 6.800 1053.160 1429.360 ;
    RECT 1055.880 6.800 1058.600 1429.360 ;
    RECT 1061.320 6.800 1064.040 1429.360 ;
    RECT 1066.760 6.800 1069.480 1429.360 ;
    RECT 1072.200 6.800 1074.920 1429.360 ;
    RECT 1077.640 6.800 1080.360 1429.360 ;
    RECT 1083.080 6.800 1085.800 1429.360 ;
    RECT 1088.520 6.800 1091.240 1429.360 ;
    RECT 1093.960 6.800 1096.680 1429.360 ;
    RECT 1099.400 6.800 1102.120 1429.360 ;
    RECT 1104.840 6.800 1107.560 1429.360 ;
    RECT 1110.280 6.800 1113.000 1429.360 ;
    RECT 1115.720 6.800 1118.440 1429.360 ;
    RECT 1121.160 6.800 1123.880 1429.360 ;
    RECT 1126.600 6.800 1129.320 1429.360 ;
    RECT 1132.040 6.800 1134.760 1429.360 ;
    RECT 1137.480 6.800 1140.200 1429.360 ;
    RECT 1142.920 6.800 1145.640 1429.360 ;
    RECT 1148.360 6.800 1151.080 1429.360 ;
    RECT 1153.800 6.800 1156.520 1429.360 ;
    RECT 1159.240 6.800 1161.960 1429.360 ;
    RECT 1164.680 6.800 1167.400 1429.360 ;
    RECT 1170.120 6.800 1172.840 1429.360 ;
    RECT 1175.560 6.800 1178.280 1429.360 ;
    RECT 1181.000 6.800 1183.720 1429.360 ;
    RECT 1186.440 6.800 1189.160 1429.360 ;
    RECT 1191.880 6.800 1194.600 1429.360 ;
    RECT 1197.320 6.800 1200.040 1429.360 ;
    RECT 1202.760 6.800 1205.480 1429.360 ;
    RECT 1208.200 6.800 1210.920 1429.360 ;
    RECT 1213.640 6.800 1216.360 1429.360 ;
    RECT 1219.080 6.800 1221.800 1429.360 ;
    RECT 1224.520 6.800 1227.240 1429.360 ;
    RECT 1229.960 6.800 1232.680 1429.360 ;
    RECT 1235.400 6.800 1238.120 1429.360 ;
    RECT 1240.840 6.800 1243.560 1429.360 ;
    RECT 1246.280 6.800 1249.000 1429.360 ;
    RECT 1251.720 6.800 1254.440 1429.360 ;
    RECT 1257.160 6.800 1259.880 1429.360 ;
    RECT 1262.600 6.800 1265.320 1429.360 ;
    RECT 1268.040 6.800 1270.760 1429.360 ;
    RECT 1273.480 6.800 1276.200 1429.360 ;
    RECT 1278.920 6.800 1281.640 1429.360 ;
    RECT 1284.360 6.800 1287.080 1429.360 ;
    RECT 1289.800 6.800 1292.520 1429.360 ;
    RECT 1295.240 6.800 1297.960 1429.360 ;
    RECT 1300.680 6.800 1303.400 1429.360 ;
    RECT 1306.120 6.800 1308.840 1429.360 ;
    RECT 1311.560 6.800 1314.280 1429.360 ;
    RECT 1317.000 6.800 1319.720 1429.360 ;
    RECT 1322.440 6.800 1325.160 1429.360 ;
    RECT 1327.880 6.800 1330.600 1429.360 ;
    RECT 1333.320 6.800 1336.040 1429.360 ;
    RECT 1338.760 6.800 1341.480 1429.360 ;
    RECT 1344.200 6.800 1346.920 1429.360 ;
    RECT 1349.640 6.800 1352.360 1429.360 ;
    RECT 1355.080 6.800 1357.800 1429.360 ;
    RECT 1360.520 6.800 1363.240 1429.360 ;
    RECT 1365.960 6.800 1368.680 1429.360 ;
    RECT 1371.400 6.800 1374.120 1429.360 ;
    RECT 1376.840 6.800 1379.560 1429.360 ;
    RECT 1382.280 6.800 1385.000 1429.360 ;
    RECT 1387.720 6.800 1390.440 1429.360 ;
    RECT 1393.160 6.800 1395.880 1429.360 ;
    RECT 1398.600 6.800 1401.320 1429.360 ;
    RECT 1404.040 6.800 1406.760 1429.360 ;
    RECT 1409.480 6.800 1412.200 1429.360 ;
    RECT 1414.920 6.800 1417.640 1429.360 ;
    RECT 1420.360 6.800 1423.080 1429.360 ;
    RECT 1425.800 6.800 1428.520 1429.360 ;
    RECT 1431.240 6.800 1433.960 1429.360 ;
    RECT 1436.680 6.800 1439.400 1429.360 ;
    RECT 1442.120 6.800 1444.840 1429.360 ;
    RECT 1447.560 6.800 1450.280 1429.360 ;
    RECT 1453.000 6.800 1455.720 1429.360 ;
    RECT 1458.440 6.800 1461.160 1429.360 ;
    RECT 1463.880 6.800 1466.600 1429.360 ;
    RECT 1469.320 6.800 1472.040 1429.360 ;
    RECT 1474.760 6.800 1477.480 1429.360 ;
    RECT 1480.200 6.800 1482.920 1429.360 ;
    RECT 1485.640 6.800 1488.360 1429.360 ;
    RECT 1491.080 6.800 1493.800 1429.360 ;
    RECT 1496.520 6.800 1499.240 1429.360 ;
    RECT 1501.960 6.800 1504.680 1429.360 ;
    RECT 1507.400 6.800 1510.120 1429.360 ;
    RECT 1512.840 6.800 1515.560 1429.360 ;
    RECT 1518.280 6.800 1521.000 1429.360 ;
    RECT 1523.720 6.800 1526.440 1429.360 ;
    RECT 1529.160 6.800 1531.880 1429.360 ;
    RECT 1534.600 6.800 1537.320 1429.360 ;
    RECT 1540.040 6.800 1542.760 1429.360 ;
    RECT 1545.480 6.800 1548.200 1429.360 ;
    RECT 1550.920 6.800 1553.640 1429.360 ;
    RECT 1556.360 6.800 1559.080 1429.360 ;
    RECT 1561.800 6.800 1564.520 1429.360 ;
    RECT 1567.240 6.800 1569.960 1429.360 ;
    RECT 1572.680 6.800 1575.400 1429.360 ;
    RECT 1578.120 6.800 1580.840 1429.360 ;
    RECT 1583.560 6.800 1586.280 1429.360 ;
    RECT 1589.000 6.800 1591.720 1429.360 ;
    RECT 1594.440 6.800 1597.160 1429.360 ;
    RECT 1599.880 6.800 1602.600 1429.360 ;
    RECT 1605.320 6.800 1608.040 1429.360 ;
    RECT 1610.760 6.800 1613.480 1429.360 ;
    RECT 1616.200 6.800 1618.920 1429.360 ;
    RECT 1621.640 6.800 1624.360 1429.360 ;
    RECT 1627.080 6.800 1629.800 1429.360 ;
    RECT 1632.520 6.800 1635.240 1429.360 ;
    RECT 1637.960 6.800 1640.680 1429.360 ;
    RECT 1643.400 6.800 1646.120 1429.360 ;
    RECT 1648.840 6.800 1651.560 1429.360 ;
    RECT 1654.280 6.800 1657.000 1429.360 ;
    RECT 1659.720 6.800 1662.440 1429.360 ;
    RECT 1665.160 6.800 1667.880 1429.360 ;
    RECT 1670.600 6.800 1673.320 1429.360 ;
    RECT 1676.040 6.800 1678.760 1429.360 ;
    RECT 1681.480 6.800 1684.200 1429.360 ;
    RECT 1686.920 6.800 1689.640 1429.360 ;
    RECT 1692.360 6.800 1695.080 1429.360 ;
    RECT 1697.800 6.800 1700.520 1429.360 ;
    RECT 1703.240 6.800 1705.960 1429.360 ;
    RECT 1708.680 6.800 1711.400 1429.360 ;
    RECT 1714.120 6.800 1716.840 1429.360 ;
    RECT 1719.560 6.800 1722.280 1429.360 ;
    RECT 1725.000 6.800 1727.720 1429.360 ;
    RECT 1730.440 6.800 1733.160 1429.360 ;
    RECT 1735.880 6.800 1738.600 1429.360 ;
    RECT 1741.320 6.800 1744.040 1429.360 ;
    RECT 1746.760 6.800 1749.480 1429.360 ;
    RECT 1752.200 6.800 1754.920 1429.360 ;
    RECT 1757.640 6.800 1760.360 1429.360 ;
    RECT 1763.080 6.800 1765.800 1429.360 ;
    RECT 1768.520 6.800 1771.240 1429.360 ;
    RECT 1773.960 6.800 1776.680 1429.360 ;
    RECT 1779.400 6.800 1782.120 1429.360 ;
    RECT 1784.840 6.800 1787.560 1429.360 ;
    RECT 1790.280 6.800 1793.000 1429.360 ;
    RECT 1795.720 6.800 1798.440 1429.360 ;
    RECT 1801.160 6.800 1803.880 1429.360 ;
    RECT 1806.600 6.800 1809.320 1429.360 ;
    RECT 1812.040 6.800 1814.760 1429.360 ;
    RECT 1817.480 6.800 1820.200 1429.360 ;
    RECT 1822.920 6.800 1825.640 1429.360 ;
    RECT 1828.360 6.800 1831.080 1429.360 ;
    RECT 1833.800 6.800 1836.520 1429.360 ;
    RECT 1839.240 6.800 1841.960 1429.360 ;
    RECT 1844.680 6.800 1847.400 1429.360 ;
    RECT 1850.120 6.800 1852.840 1429.360 ;
    RECT 1855.560 6.800 1858.280 1429.360 ;
    RECT 1861.000 6.800 1863.720 1429.360 ;
    RECT 1866.440 6.800 1869.160 1429.360 ;
    RECT 1871.880 6.800 1874.600 1429.360 ;
    RECT 1877.320 6.800 1880.040 1429.360 ;
    RECT 1882.760 6.800 1885.480 1429.360 ;
    RECT 1888.200 6.800 1890.920 1429.360 ;
    RECT 1893.640 6.800 1896.360 1429.360 ;
    RECT 1899.080 6.800 1901.800 1429.360 ;
    RECT 1904.520 6.800 1907.240 1429.360 ;
    RECT 1909.960 6.800 1912.680 1429.360 ;
    RECT 1915.400 6.800 1918.120 1429.360 ;
    RECT 1920.840 6.800 1923.560 1429.360 ;
    RECT 1926.280 6.800 1929.000 1429.360 ;
    RECT 1931.720 6.800 1934.440 1429.360 ;
    RECT 1937.160 6.800 1939.880 1429.360 ;
    RECT 1942.600 6.800 1945.320 1429.360 ;
    RECT 1948.040 6.800 1950.760 1429.360 ;
    RECT 1953.480 6.800 1956.200 1429.360 ;
    RECT 1958.920 6.800 1961.640 1429.360 ;
    RECT 1964.360 6.800 1967.080 1429.360 ;
    RECT 1969.800 6.800 1972.520 1429.360 ;
    RECT 1975.240 6.800 1977.960 1429.360 ;
    RECT 1980.680 6.800 1983.400 1429.360 ;
    RECT 1986.120 6.800 1988.840 1429.360 ;
    RECT 1991.560 6.800 1994.280 1429.360 ;
    RECT 1997.000 6.800 1999.720 1429.360 ;
    RECT 2002.440 6.800 2005.160 1429.360 ;
    RECT 2007.880 6.800 2010.600 1429.360 ;
    RECT 2013.320 6.800 2016.040 1429.360 ;
    RECT 2018.760 6.800 2021.480 1429.360 ;
    RECT 2024.200 6.800 2026.920 1429.360 ;
    RECT 2029.640 6.800 2032.360 1429.360 ;
    RECT 2035.080 6.800 2037.800 1429.360 ;
    RECT 2040.520 6.800 2043.240 1429.360 ;
    RECT 2045.960 6.800 2048.680 1429.360 ;
    RECT 2051.400 6.800 2054.120 1429.360 ;
    RECT 2056.840 6.800 2059.560 1429.360 ;
    RECT 2062.280 6.800 2065.000 1429.360 ;
    RECT 2067.720 6.800 2070.440 1429.360 ;
    RECT 2073.160 6.800 2075.880 1429.360 ;
    RECT 2078.600 6.800 2081.320 1429.360 ;
    RECT 2084.040 6.800 2086.760 1429.360 ;
    RECT 2089.480 6.800 2092.200 1429.360 ;
    RECT 2094.920 6.800 2097.640 1429.360 ;
    RECT 2100.360 6.800 2103.080 1429.360 ;
    RECT 2105.800 6.800 2108.520 1429.360 ;
    RECT 2111.240 6.800 2113.960 1429.360 ;
    RECT 2116.680 6.800 2119.400 1429.360 ;
    RECT 2122.120 6.800 2124.840 1429.360 ;
    RECT 2127.560 6.800 2130.280 1429.360 ;
    RECT 2133.000 6.800 2135.720 1429.360 ;
    RECT 2138.440 6.800 2141.160 1429.360 ;
    RECT 2143.880 6.800 2146.600 1429.360 ;
    RECT 2149.320 6.800 2152.040 1429.360 ;
    RECT 2154.760 6.800 2157.480 1429.360 ;
    RECT 2160.200 6.800 2162.920 1429.360 ;
    RECT 2165.640 6.800 2168.360 1429.360 ;
    RECT 2171.080 6.800 2173.800 1429.360 ;
    RECT 2176.520 6.800 2179.240 1429.360 ;
    RECT 2181.960 6.800 2184.680 1429.360 ;
    RECT 2187.400 6.800 2190.120 1429.360 ;
    RECT 2192.840 6.800 2195.560 1429.360 ;
    RECT 2198.280 6.800 2201.000 1429.360 ;
    RECT 2203.720 6.800 2206.440 1429.360 ;
    RECT 2209.160 6.800 2211.880 1429.360 ;
    RECT 2214.600 6.800 2217.320 1429.360 ;
    RECT 2220.040 6.800 2222.760 1429.360 ;
    RECT 2225.480 6.800 2228.200 1429.360 ;
    RECT 2230.920 6.800 2233.640 1429.360 ;
    RECT 2236.360 6.800 2239.080 1429.360 ;
    RECT 2241.800 6.800 2244.520 1429.360 ;
    RECT 2247.240 6.800 2249.960 1429.360 ;
    RECT 2252.680 6.800 2255.400 1429.360 ;
    RECT 2258.120 6.800 2260.840 1429.360 ;
    RECT 2263.560 6.800 2266.280 1429.360 ;
    RECT 2269.000 6.800 2271.720 1429.360 ;
    RECT 2274.440 6.800 2277.160 1429.360 ;
    RECT 2279.880 6.800 2282.600 1429.360 ;
    RECT 2285.320 6.800 2288.040 1429.360 ;
    RECT 2290.760 6.800 2293.480 1429.360 ;
    RECT 2296.200 6.800 2298.920 1429.360 ;
    RECT 2301.640 6.800 2304.360 1429.360 ;
    RECT 2307.080 6.800 2309.800 1429.360 ;
    RECT 2312.520 6.800 2315.240 1429.360 ;
    RECT 2317.960 6.800 2320.680 1429.360 ;
    RECT 2323.400 6.800 2326.120 1429.360 ;
    RECT 2328.840 6.800 2331.560 1429.360 ;
    RECT 2334.280 6.800 2337.000 1429.360 ;
    RECT 2339.720 6.800 2342.440 1429.360 ;
    RECT 2345.160 6.800 2347.880 1429.360 ;
    RECT 2350.600 6.800 2353.320 1429.360 ;
    RECT 2356.040 6.800 2358.760 1429.360 ;
    RECT 2361.480 6.800 2364.200 1429.360 ;
    RECT 2366.920 6.800 2369.640 1429.360 ;
    RECT 2372.360 6.800 2375.080 1429.360 ;
    RECT 2377.800 6.800 2380.520 1429.360 ;
    RECT 2383.240 6.800 2385.960 1429.360 ;
    RECT 2388.680 6.800 2391.400 1429.360 ;
    RECT 2394.120 6.800 2396.840 1429.360 ;
    RECT 2399.560 6.800 2402.280 1429.360 ;
    RECT 2405.000 6.800 2407.720 1429.360 ;
    RECT 2410.440 6.800 2413.160 1429.360 ;
    RECT 2415.880 6.800 2418.600 1429.360 ;
    RECT 2421.320 6.800 2424.040 1429.360 ;
    RECT 2426.760 6.800 2429.480 1429.360 ;
    RECT 2432.200 6.800 2434.920 1429.360 ;
    RECT 2437.640 6.800 2440.360 1429.360 ;
    RECT 2443.080 6.800 2445.800 1429.360 ;
    RECT 2448.520 6.800 2451.240 1429.360 ;
    RECT 2453.960 6.800 2456.680 1429.360 ;
    RECT 2459.400 6.800 2462.120 1429.360 ;
    RECT 2464.840 6.800 2467.560 1429.360 ;
    RECT 2470.280 6.800 2473.000 1429.360 ;
    RECT 2475.720 6.800 2478.440 1429.360 ;
    RECT 2481.160 6.800 2483.880 1429.360 ;
    RECT 2486.600 6.800 2489.320 1429.360 ;
    RECT 2492.040 6.800 2494.760 1429.360 ;
    RECT 2497.480 6.800 2500.200 1429.360 ;
    RECT 2502.920 6.800 2505.640 1429.360 ;
    RECT 2508.360 6.800 2511.080 1429.360 ;
    RECT 2513.800 6.800 2516.520 1429.360 ;
    RECT 2519.240 6.800 2521.960 1429.360 ;
    RECT 2524.680 6.800 2527.400 1429.360 ;
    RECT 2530.120 6.800 2532.840 1429.360 ;
    RECT 2535.560 6.800 2538.280 1429.360 ;
    RECT 2541.000 6.800 2543.720 1429.360 ;
    RECT 2546.440 6.800 2549.160 1429.360 ;
    RECT 2551.880 6.800 2554.600 1429.360 ;
    RECT 2557.320 6.800 2560.040 1429.360 ;
    RECT 2562.760 6.800 2565.480 1429.360 ;
    RECT 2568.200 6.800 2570.920 1429.360 ;
    RECT 2573.640 6.800 2576.360 1429.360 ;
    RECT 2579.080 6.800 2581.800 1429.360 ;
    RECT 2584.520 6.800 2587.240 1429.360 ;
    RECT 2589.960 6.800 2592.680 1429.360 ;
    RECT 2595.400 6.800 2598.120 1429.360 ;
    RECT 2600.840 6.800 2603.560 1429.360 ;
    RECT 2606.280 6.800 2609.000 1429.360 ;
    RECT 2611.720 6.800 2614.440 1429.360 ;
    RECT 2617.160 6.800 2619.880 1429.360 ;
    RECT 2622.600 6.800 2625.320 1429.360 ;
    RECT 2628.040 6.800 2630.760 1429.360 ;
    RECT 2633.480 6.800 2636.200 1429.360 ;
    RECT 2638.920 6.800 2641.640 1429.360 ;
    RECT 2644.360 6.800 2647.080 1429.360 ;
    RECT 2649.800 6.800 2652.520 1429.360 ;
    RECT 2655.240 6.800 2657.960 1429.360 ;
    RECT 2660.680 6.800 2663.400 1429.360 ;
    RECT 2666.120 6.800 2668.840 1429.360 ;
    RECT 2671.560 6.800 2674.280 1429.360 ;
    RECT 2677.000 6.800 2679.720 1429.360 ;
    RECT 2682.440 6.800 2685.160 1429.360 ;
    RECT 2687.880 6.800 2690.600 1429.360 ;
    RECT 2693.320 6.800 2696.040 1429.360 ;
    RECT 2698.760 6.800 2701.480 1429.360 ;
    RECT 2704.200 6.800 2706.920 1429.360 ;
    RECT 2709.640 6.800 2712.360 1429.360 ;
    RECT 2715.080 6.800 2717.800 1429.360 ;
    RECT 2720.520 6.800 2723.240 1429.360 ;
    RECT 2725.960 6.800 2728.680 1429.360 ;
    RECT 2731.400 6.800 2734.120 1429.360 ;
    RECT 2736.840 6.800 2739.560 1429.360 ;
    RECT 2742.280 6.800 2745.000 1429.360 ;
    RECT 2747.720 6.800 2750.440 1429.360 ;
    RECT 2753.160 6.800 2755.880 1429.360 ;
    RECT 2758.600 6.800 2761.320 1429.360 ;
    RECT 2764.040 6.800 2766.760 1429.360 ;
    RECT 2769.480 6.800 2772.200 1429.360 ;
    RECT 2774.920 6.800 2777.640 1429.360 ;
    RECT 2780.360 6.800 2783.080 1429.360 ;
    RECT 2785.800 6.800 2788.520 1429.360 ;
    RECT 2791.240 6.800 2793.960 1429.360 ;
    RECT 2796.680 6.800 2799.400 1429.360 ;
    RECT 2802.120 6.800 2804.840 1429.360 ;
    RECT 2807.560 6.800 2810.280 1429.360 ;
    RECT 2813.000 6.800 2815.720 1429.360 ;
    RECT 2818.440 6.800 2821.160 1429.360 ;
    RECT 2823.880 6.800 2826.600 1429.360 ;
    RECT 2829.320 6.800 2832.040 1429.360 ;
    RECT 2834.760 6.800 2837.480 1429.360 ;
    RECT 2840.200 6.800 2842.920 1429.360 ;
    RECT 2845.640 6.800 2848.360 1429.360 ;
    RECT 2851.080 6.800 2853.800 1429.360 ;
    RECT 2856.520 6.800 2859.240 1429.360 ;
    RECT 2861.960 6.800 2864.680 1429.360 ;
    RECT 2867.400 6.800 2870.120 1429.360 ;
    RECT 2872.840 6.800 2875.560 1429.360 ;
    RECT 2878.280 6.800 2881.000 1429.360 ;
    RECT 2883.720 6.800 2886.440 1429.360 ;
    RECT 2889.160 6.800 2891.880 1429.360 ;
    RECT 2894.600 6.800 2897.320 1429.360 ;
    RECT 2900.040 6.800 2902.760 1429.360 ;
    RECT 2905.480 6.800 2908.200 1429.360 ;
    RECT 2910.920 6.800 2913.640 1429.360 ;
    RECT 2916.360 6.800 2919.080 1429.360 ;
    RECT 2921.800 6.800 2924.520 1429.360 ;
    RECT 2927.240 6.800 2929.960 1429.360 ;
    RECT 2932.680 6.800 2935.400 1429.360 ;
    RECT 2938.120 6.800 2940.840 1429.360 ;
    RECT 2943.560 6.800 2946.280 1429.360 ;
    RECT 2949.000 6.800 2951.720 1429.360 ;
    RECT 2954.440 6.800 2957.160 1429.360 ;
    RECT 2959.880 6.800 2962.600 1429.360 ;
    RECT 2965.320 6.800 2968.040 1429.360 ;
    RECT 2970.760 6.800 2973.480 1429.360 ;
    RECT 2976.200 6.800 2978.920 1429.360 ;
    RECT 2981.640 6.800 2984.360 1429.360 ;
    RECT 2987.080 6.800 2989.800 1429.360 ;
    RECT 2992.520 6.800 2995.240 1429.360 ;
    RECT 2997.960 6.800 3000.680 1429.360 ;
    RECT 3003.400 6.800 3006.120 1429.360 ;
    RECT 3008.840 6.800 3011.560 1429.360 ;
    RECT 3014.280 6.800 3017.000 1429.360 ;
    RECT 3019.720 6.800 3022.440 1429.360 ;
    RECT 3025.160 6.800 3027.880 1429.360 ;
    RECT 3030.600 6.800 3033.320 1429.360 ;
    RECT 3036.040 6.800 3038.760 1429.360 ;
    RECT 3041.480 6.800 3044.200 1429.360 ;
    RECT 3046.920 6.800 3049.640 1429.360 ;
    RECT 3052.360 6.800 3055.080 1429.360 ;
    RECT 3057.800 6.800 3060.520 1429.360 ;
    RECT 3063.240 6.800 3065.960 1429.360 ;
    RECT 3068.680 6.800 3071.400 1429.360 ;
    RECT 3074.120 6.800 3076.840 1429.360 ;
    RECT 3079.560 6.800 3082.280 1429.360 ;
    RECT 3085.000 6.800 3087.720 1429.360 ;
    RECT 3090.440 6.800 3093.160 1429.360 ;
    RECT 3095.880 6.800 3098.600 1429.360 ;
    RECT 3101.320 6.800 3104.040 1429.360 ;
    RECT 3106.760 6.800 3109.480 1429.360 ;
    RECT 3112.200 6.800 3114.920 1429.360 ;
    RECT 3117.640 6.800 3120.360 1429.360 ;
    RECT 3123.080 6.800 3125.800 1429.360 ;
    RECT 3128.520 6.800 3131.240 1429.360 ;
    RECT 3133.960 6.800 3136.680 1429.360 ;
    RECT 3139.400 6.800 3142.120 1429.360 ;
    RECT 3144.840 6.800 3147.560 1429.360 ;
    RECT 3150.280 6.800 3153.000 1429.360 ;
    RECT 3155.720 6.800 3158.440 1429.360 ;
    RECT 3161.160 6.800 3163.880 1429.360 ;
    RECT 3166.600 6.800 3169.320 1429.360 ;
    RECT 3172.040 6.800 3174.760 1429.360 ;
    RECT 3177.480 6.800 3180.200 1429.360 ;
    RECT 3182.920 6.800 3185.640 1429.360 ;
    RECT 3188.360 6.800 3191.080 1429.360 ;
    RECT 3193.800 6.800 3196.520 1429.360 ;
    RECT 3199.240 6.800 3201.960 1429.360 ;
    RECT 3204.680 6.800 3207.400 1429.360 ;
    RECT 3210.120 6.800 3212.840 1429.360 ;
    RECT 3215.560 6.800 3218.280 1429.360 ;
    RECT 3221.000 6.800 3223.720 1429.360 ;
    RECT 3226.440 6.800 3229.160 1429.360 ;
    RECT 3231.880 6.800 3234.600 1429.360 ;
    RECT 3237.320 6.800 3240.040 1429.360 ;
    RECT 3242.760 6.800 3245.480 1429.360 ;
    RECT 3248.200 6.800 3250.920 1429.360 ;
    RECT 3253.640 6.800 3256.360 1429.360 ;
    RECT 3259.080 6.800 3261.800 1429.360 ;
    RECT 3264.520 6.800 3267.240 1429.360 ;
    RECT 3269.960 6.800 3272.680 1429.360 ;
    RECT 3275.400 6.800 3278.120 1429.360 ;
    RECT 3280.840 6.800 3283.560 1429.360 ;
    RECT 3286.280 6.800 3289.000 1429.360 ;
    RECT 3291.720 6.800 3294.440 1429.360 ;
    RECT 3297.160 6.800 3299.880 1429.360 ;
    RECT 3302.600 6.800 3305.320 1429.360 ;
    RECT 3308.040 6.800 3310.760 1429.360 ;
    RECT 3313.480 6.800 3316.200 1429.360 ;
    RECT 3318.920 6.800 3321.640 1429.360 ;
    RECT 3324.360 6.800 3327.080 1429.360 ;
    RECT 3329.800 6.800 3332.520 1429.360 ;
    RECT 3335.240 6.800 3337.960 1429.360 ;
    RECT 3340.680 6.800 3343.400 1429.360 ;
    RECT 3346.120 6.800 3348.840 1429.360 ;
    RECT 3351.560 6.800 3354.280 1429.360 ;
    RECT 3357.000 6.800 3359.720 1429.360 ;
    RECT 3362.440 6.800 3365.160 1429.360 ;
    RECT 3367.880 6.800 3370.600 1429.360 ;
    RECT 3373.320 6.800 3376.040 1429.360 ;
    RECT 3378.760 6.800 3381.480 1429.360 ;
    RECT 3384.200 6.800 3386.920 1429.360 ;
    RECT 3389.640 6.800 3392.360 1429.360 ;
    RECT 3395.080 6.800 3397.800 1429.360 ;
    RECT 3400.520 6.800 3403.240 1429.360 ;
    RECT 3405.960 6.800 3408.680 1429.360 ;
    RECT 3411.400 6.800 3414.120 1429.360 ;
    RECT 3416.840 6.800 3419.560 1429.360 ;
    RECT 3422.280 6.800 3425.000 1429.360 ;
    RECT 3427.720 6.800 3430.440 1429.360 ;
    RECT 3433.160 6.800 3435.880 1429.360 ;
    RECT 3438.600 6.800 3441.320 1429.360 ;
    RECT 3444.040 6.800 3446.760 1429.360 ;
    RECT 3449.480 6.800 3452.200 1429.360 ;
    RECT 3454.920 6.800 3457.640 1429.360 ;
    RECT 3460.360 6.800 3463.080 1429.360 ;
    RECT 3465.800 6.800 3468.520 1429.360 ;
    RECT 3471.240 6.800 3473.960 1429.360 ;
    RECT 3476.680 6.800 3479.400 1429.360 ;
    RECT 3482.120 6.800 3484.840 1429.360 ;
    RECT 3487.560 6.800 3490.280 1429.360 ;
    RECT 3493.000 6.800 3495.720 1429.360 ;
    RECT 3498.440 6.800 3501.160 1429.360 ;
    RECT 3503.880 6.800 3506.600 1429.360 ;
    RECT 3509.320 6.800 3512.040 1429.360 ;
    RECT 3514.760 6.800 3517.480 1429.360 ;
    RECT 3520.200 6.800 3522.920 1429.360 ;
    RECT 3525.640 6.800 3528.360 1429.360 ;
    RECT 3531.080 6.800 3533.800 1429.360 ;
    RECT 3536.520 6.800 3539.240 1429.360 ;
    RECT 3541.960 6.800 3544.680 1429.360 ;
    RECT 3547.400 6.800 3550.120 1429.360 ;
    RECT 3552.840 6.800 3555.560 1429.360 ;
    RECT 3558.280 6.800 3561.000 1429.360 ;
    RECT 3563.720 6.800 3566.440 1429.360 ;
    RECT 3569.160 6.800 3571.880 1429.360 ;
    RECT 3574.600 6.800 3577.320 1429.360 ;
    RECT 3580.040 6.800 3582.760 1429.360 ;
    RECT 3585.480 6.800 3588.200 1429.360 ;
    RECT 3590.920 6.800 3593.640 1429.360 ;
    RECT 3596.360 6.800 3599.080 1429.360 ;
    RECT 3601.800 6.800 3604.520 1429.360 ;
    RECT 3607.240 6.800 3609.960 1429.360 ;
    RECT 3612.680 6.800 3615.400 1429.360 ;
    RECT 3618.120 6.800 3620.840 1429.360 ;
    RECT 3623.560 6.800 3626.280 1429.360 ;
    RECT 3629.000 6.800 3631.720 1429.360 ;
    RECT 3634.440 6.800 3637.160 1429.360 ;
    RECT 3639.880 6.800 3642.600 1429.360 ;
    RECT 3645.320 6.800 3648.040 1429.360 ;
    RECT 3650.760 6.800 3653.480 1429.360 ;
    RECT 3656.200 6.800 3658.920 1429.360 ;
    RECT 3661.640 6.800 3664.360 1429.360 ;
    RECT 3667.080 6.800 3669.800 1429.360 ;
    RECT 3672.520 6.800 3675.240 1429.360 ;
    RECT 3677.960 6.800 3680.680 1429.360 ;
    RECT 3683.400 6.800 3686.120 1429.360 ;
    RECT 3688.840 6.800 3691.560 1429.360 ;
    RECT 3694.280 6.800 3697.000 1429.360 ;
    RECT 3699.720 6.800 3702.440 1429.360 ;
    RECT 3705.160 6.800 3707.880 1429.360 ;
    RECT 3710.600 6.800 3713.320 1429.360 ;
    RECT 3716.040 6.800 3718.760 1429.360 ;
    RECT 3721.480 6.800 3724.200 1429.360 ;
    RECT 3726.920 6.800 3729.640 1429.360 ;
    RECT 3732.360 6.800 3735.080 1429.360 ;
    RECT 3737.800 6.800 3740.520 1429.360 ;
    RECT 3743.240 6.800 3745.960 1429.360 ;
    RECT 3748.680 6.800 3751.400 1429.360 ;
    RECT 3754.120 6.800 3756.840 1429.360 ;
    RECT 3759.560 6.800 3762.280 1429.360 ;
    RECT 3765.000 6.800 3767.720 1429.360 ;
    RECT 3770.440 6.800 3773.160 1429.360 ;
    RECT 3775.880 6.800 3778.600 1429.360 ;
    RECT 3781.320 6.800 3784.040 1429.360 ;
    RECT 3786.760 6.800 3789.480 1429.360 ;
    RECT 3792.200 6.800 3794.920 1429.360 ;
    RECT 3797.640 6.800 3800.360 1429.360 ;
    RECT 3803.080 6.800 3805.800 1429.360 ;
    RECT 3808.520 6.800 3811.240 1429.360 ;
    RECT 3813.960 6.800 3816.680 1429.360 ;
    RECT 3819.400 6.800 3822.120 1429.360 ;
    RECT 3824.840 6.800 3827.560 1429.360 ;
    RECT 3830.280 6.800 3833.000 1429.360 ;
    RECT 3835.720 6.800 3838.440 1429.360 ;
    RECT 3841.160 6.800 3843.880 1429.360 ;
    RECT 3846.600 6.800 3849.320 1429.360 ;
    RECT 3852.040 6.800 3854.760 1429.360 ;
    RECT 3857.480 6.800 3860.200 1429.360 ;
    RECT 3862.920 6.800 3865.640 1429.360 ;
    RECT 3868.360 6.800 3871.080 1429.360 ;
    RECT 3873.800 6.800 3876.520 1429.360 ;
    RECT 3879.240 6.800 3881.960 1429.360 ;
    RECT 3884.680 6.800 3887.400 1429.360 ;
    RECT 3890.120 6.800 3892.840 1429.360 ;
    RECT 3895.560 6.800 3898.280 1429.360 ;
    RECT 3901.000 6.800 3903.720 1429.360 ;
    RECT 3906.440 6.800 3909.160 1429.360 ;
    RECT 3911.880 6.800 3914.600 1429.360 ;
    RECT 3917.320 6.800 3920.040 1429.360 ;
    RECT 3922.760 6.800 3925.480 1429.360 ;
    RECT 3928.200 6.800 3930.920 1429.360 ;
    RECT 3933.640 6.800 3936.360 1429.360 ;
    RECT 3939.080 6.800 3941.800 1429.360 ;
    RECT 3944.520 6.800 3947.240 1429.360 ;
    RECT 3949.960 6.800 3952.680 1429.360 ;
    RECT 3955.400 6.800 3958.120 1429.360 ;
    RECT 3960.840 6.800 3963.560 1429.360 ;
    RECT 3966.280 6.800 3969.000 1429.360 ;
    RECT 3971.720 6.800 3974.440 1429.360 ;
    RECT 3977.160 6.800 3979.880 1429.360 ;
    RECT 3982.600 6.800 3985.320 1429.360 ;
    RECT 3988.040 6.800 3990.760 1429.360 ;
    RECT 3993.480 6.800 3996.200 1429.360 ;
    RECT 3998.920 6.800 4001.640 1429.360 ;
    RECT 4004.360 6.800 4007.080 1429.360 ;
    RECT 4009.800 6.800 4012.520 1429.360 ;
    RECT 4015.240 6.800 4017.960 1429.360 ;
    RECT 4020.680 6.800 4023.400 1429.360 ;
    RECT 4026.120 6.800 4028.840 1429.360 ;
    RECT 4031.560 6.800 4034.280 1429.360 ;
    RECT 4037.000 6.800 4039.720 1429.360 ;
    RECT 4042.440 6.800 4045.160 1429.360 ;
    RECT 4047.880 6.800 4050.600 1429.360 ;
    RECT 4053.320 6.800 4056.040 1429.360 ;
    RECT 4058.760 6.800 4061.480 1429.360 ;
    RECT 4064.200 6.800 4066.920 1429.360 ;
    RECT 4069.640 6.800 4072.360 1429.360 ;
    RECT 4075.080 6.800 4077.800 1429.360 ;
    RECT 4080.520 6.800 4083.240 1429.360 ;
    RECT 4085.960 6.800 4088.680 1429.360 ;
    RECT 4091.400 6.800 4094.120 1429.360 ;
    RECT 4096.840 6.800 4099.560 1429.360 ;
    RECT 4102.280 6.800 4105.000 1429.360 ;
    RECT 4107.720 6.800 4110.440 1429.360 ;
    RECT 4113.160 6.800 4115.880 1429.360 ;
    RECT 4118.600 6.800 4121.320 1429.360 ;
    RECT 4124.040 6.800 4126.760 1429.360 ;
    RECT 4129.480 6.800 4132.200 1429.360 ;
    RECT 4134.920 6.800 4137.640 1429.360 ;
    RECT 4140.360 6.800 4143.080 1429.360 ;
    RECT 4145.800 6.800 4148.520 1429.360 ;
    RECT 4151.240 6.800 4153.960 1429.360 ;
    RECT 4156.680 6.800 4159.400 1429.360 ;
    RECT 4162.120 6.800 4164.840 1429.360 ;
    RECT 4167.560 6.800 4170.280 1429.360 ;
    RECT 4173.000 6.800 4175.720 1429.360 ;
    RECT 4178.440 6.800 4181.160 1429.360 ;
    RECT 4183.880 6.800 4186.600 1429.360 ;
    RECT 4189.320 6.800 4192.040 1429.360 ;
    RECT 4194.760 6.800 4197.480 1429.360 ;
    RECT 4200.200 6.800 4202.920 1429.360 ;
    RECT 4205.640 6.800 4208.360 1429.360 ;
    RECT 4211.080 6.800 4213.800 1429.360 ;
    RECT 4216.520 6.800 4219.240 1429.360 ;
    RECT 4221.960 6.800 4224.680 1429.360 ;
    RECT 4227.400 6.800 4230.120 1429.360 ;
    RECT 4232.840 6.800 4235.560 1429.360 ;
    RECT 4238.280 6.800 4241.000 1429.360 ;
    RECT 4243.720 6.800 4246.440 1429.360 ;
    RECT 4249.160 6.800 4251.880 1429.360 ;
    RECT 4254.600 6.800 4257.320 1429.360 ;
    RECT 4260.040 6.800 4262.760 1429.360 ;
    RECT 4265.480 6.800 4268.200 1429.360 ;
    RECT 4270.920 6.800 4273.640 1429.360 ;
    RECT 4276.360 6.800 4279.080 1429.360 ;
    RECT 4281.800 6.800 4284.520 1429.360 ;
    RECT 4287.240 6.800 4289.960 1429.360 ;
    RECT 4292.680 6.800 4295.400 1429.360 ;
    RECT 4298.120 6.800 4300.840 1429.360 ;
    RECT 4303.560 6.800 4306.280 1429.360 ;
    RECT 4309.000 6.800 4311.720 1429.360 ;
    RECT 4314.440 6.800 4317.160 1429.360 ;
    RECT 4319.880 6.800 4322.600 1429.360 ;
    RECT 4325.320 6.800 4328.040 1429.360 ;
    RECT 4330.760 6.800 4333.480 1429.360 ;
    RECT 4336.200 6.800 4338.920 1429.360 ;
    RECT 4341.640 6.800 4344.360 1429.360 ;
    RECT 4347.080 6.800 4349.800 1429.360 ;
    RECT 4352.520 6.800 4355.240 1429.360 ;
    RECT 4357.960 6.800 4360.680 1429.360 ;
    RECT 4363.400 6.800 4366.120 1429.360 ;
    RECT 4368.840 6.800 4371.560 1429.360 ;
    RECT 4374.280 6.800 4377.000 1429.360 ;
    RECT 4379.720 6.800 4382.440 1429.360 ;
    RECT 4385.160 6.800 4387.880 1429.360 ;
    RECT 4390.600 6.800 4393.320 1429.360 ;
    RECT 4396.040 6.800 4398.760 1429.360 ;
    RECT 4401.480 6.800 4404.200 1429.360 ;
    RECT 4406.920 6.800 4409.640 1429.360 ;
    RECT 4412.360 6.800 4415.080 1429.360 ;
    RECT 4417.800 6.800 4420.520 1429.360 ;
    RECT 4423.240 6.800 4425.960 1429.360 ;
    RECT 4428.680 6.800 4431.400 1429.360 ;
    RECT 4434.120 6.800 4436.840 1429.360 ;
    RECT 4439.560 6.800 4442.280 1429.360 ;
    RECT 4445.000 6.800 4447.720 1429.360 ;
    RECT 4450.440 6.800 4453.160 1429.360 ;
    RECT 4455.880 6.800 4458.600 1429.360 ;
    RECT 4461.320 6.800 4464.040 1429.360 ;
    RECT 4466.760 6.800 4469.480 1429.360 ;
    RECT 4472.200 6.800 4474.920 1429.360 ;
    RECT 4477.640 6.800 4480.360 1429.360 ;
    RECT 4483.080 6.800 4485.800 1429.360 ;
    RECT 4488.520 6.800 4491.240 1429.360 ;
    RECT 4493.960 6.800 4496.680 1429.360 ;
    RECT 4499.400 6.800 4502.120 1429.360 ;
    RECT 4504.840 6.800 4507.560 1429.360 ;
    RECT 4510.280 6.800 4513.000 1429.360 ;
    RECT 4515.720 6.800 4518.440 1429.360 ;
    RECT 4521.160 6.800 4523.880 1429.360 ;
    RECT 4526.600 6.800 4529.320 1429.360 ;
    RECT 4532.040 6.800 4534.760 1429.360 ;
    RECT 4537.480 6.800 4540.200 1429.360 ;
    RECT 4542.920 6.800 4545.640 1429.360 ;
    RECT 4548.360 6.800 4551.080 1429.360 ;
    RECT 4553.800 6.800 4556.520 1429.360 ;
    RECT 4559.240 6.800 4561.960 1429.360 ;
    RECT 4564.680 6.800 4567.400 1429.360 ;
    RECT 4570.120 6.800 4572.840 1429.360 ;
    RECT 4575.560 6.800 4578.280 1429.360 ;
    RECT 4581.000 6.800 4583.720 1429.360 ;
    RECT 4586.440 6.800 4589.160 1429.360 ;
    RECT 4591.880 6.800 4594.600 1429.360 ;
    RECT 4597.320 6.800 4600.040 1429.360 ;
    RECT 4602.760 6.800 4605.480 1429.360 ;
    RECT 4608.200 6.800 4610.920 1429.360 ;
    RECT 4613.640 6.800 4616.360 1429.360 ;
    RECT 4619.080 6.800 4621.800 1429.360 ;
    RECT 4624.520 6.800 4627.240 1429.360 ;
    RECT 4629.960 6.800 4632.680 1429.360 ;
    RECT 4635.400 6.800 4638.120 1429.360 ;
    RECT 4640.840 6.800 4643.560 1429.360 ;
    RECT 4646.280 6.800 4649.000 1429.360 ;
    RECT 4651.720 6.800 4654.440 1429.360 ;
    RECT 4657.160 6.800 4659.880 1429.360 ;
    RECT 4662.600 6.800 4665.320 1429.360 ;
    RECT 4668.040 6.800 4670.760 1429.360 ;
    RECT 4673.480 6.800 4676.200 1429.360 ;
    RECT 4678.920 6.800 4681.640 1429.360 ;
    RECT 4684.360 6.800 4687.080 1429.360 ;
    RECT 4689.800 6.800 4692.520 1429.360 ;
    RECT 4695.240 6.800 4697.960 1429.360 ;
    RECT 4700.680 6.800 4703.400 1429.360 ;
    RECT 4706.120 6.800 4708.840 1429.360 ;
    RECT 4711.560 6.800 4714.280 1429.360 ;
    RECT 4717.000 6.800 4719.720 1429.360 ;
    RECT 4722.440 6.800 4725.160 1429.360 ;
    RECT 4727.880 6.800 4730.600 1429.360 ;
    RECT 4733.320 6.800 4736.040 1429.360 ;
    RECT 4738.760 6.800 4741.480 1429.360 ;
    RECT 4744.200 6.800 4746.920 1429.360 ;
    RECT 4749.640 6.800 4752.360 1429.360 ;
    RECT 4755.080 6.800 4757.800 1429.360 ;
    RECT 4760.520 6.800 4763.240 1429.360 ;
    RECT 4765.960 6.800 4768.680 1429.360 ;
    RECT 4771.400 6.800 4774.120 1429.360 ;
    RECT 4776.840 6.800 4779.560 1429.360 ;
    RECT 4782.280 6.800 4785.000 1429.360 ;
    RECT 4787.720 6.800 4790.440 1429.360 ;
    RECT 4793.160 6.800 4795.880 1429.360 ;
    RECT 4798.600 6.800 4801.320 1429.360 ;
    RECT 4804.040 6.800 4806.760 1429.360 ;
    RECT 4809.480 6.800 4812.200 1429.360 ;
    RECT 4814.920 6.800 4817.640 1429.360 ;
    RECT 4820.360 6.800 4823.080 1429.360 ;
    RECT 4825.800 6.800 4828.520 1429.360 ;
    RECT 4831.240 6.800 4833.960 1429.360 ;
    RECT 4836.680 6.800 4839.400 1429.360 ;
    RECT 4842.120 6.800 4844.840 1429.360 ;
    RECT 4847.560 6.800 4850.280 1429.360 ;
    RECT 4853.000 6.800 4855.720 1429.360 ;
    RECT 4858.440 6.800 4861.160 1429.360 ;
    RECT 4863.880 6.800 4866.600 1429.360 ;
    RECT 4869.320 6.800 4872.040 1429.360 ;
    RECT 4874.760 6.800 4877.480 1429.360 ;
    RECT 4880.200 6.800 4882.920 1429.360 ;
    RECT 4885.640 6.800 4888.360 1429.360 ;
    RECT 4891.080 6.800 4893.800 1429.360 ;
    RECT 4896.520 6.800 4899.240 1429.360 ;
    RECT 4901.960 6.800 4904.680 1429.360 ;
    RECT 4907.400 6.800 4910.120 1429.360 ;
    RECT 4912.840 6.800 4915.560 1429.360 ;
    RECT 4918.280 6.800 4921.000 1429.360 ;
    RECT 4923.720 6.800 4926.440 1429.360 ;
    RECT 4929.160 6.800 4931.880 1429.360 ;
    RECT 4934.600 6.800 4937.320 1429.360 ;
    RECT 4940.040 6.800 4942.760 1429.360 ;
    RECT 4945.480 6.800 4948.200 1429.360 ;
    RECT 4950.920 6.800 4953.640 1429.360 ;
    RECT 4956.360 6.800 4959.080 1429.360 ;
    RECT 4961.800 6.800 4964.520 1429.360 ;
    RECT 4967.240 6.800 4969.960 1429.360 ;
    RECT 4972.680 6.800 4975.400 1429.360 ;
    RECT 4978.120 6.800 4980.840 1429.360 ;
    RECT 4983.560 6.800 4986.280 1429.360 ;
    RECT 4989.000 6.800 4991.720 1429.360 ;
    RECT 4994.440 6.800 4997.160 1429.360 ;
    RECT 4999.880 6.800 5002.600 1429.360 ;
    RECT 5005.320 6.800 5008.040 1429.360 ;
    RECT 5010.760 6.800 5013.480 1429.360 ;
    RECT 5016.200 6.800 5018.920 1429.360 ;
    RECT 5021.640 6.800 5024.360 1429.360 ;
    RECT 5027.080 6.800 5029.800 1429.360 ;
    RECT 5032.520 6.800 5035.240 1429.360 ;
    RECT 5037.960 6.800 5040.680 1429.360 ;
    RECT 5043.400 6.800 5046.120 1429.360 ;
    RECT 5048.840 6.800 5051.560 1429.360 ;
    RECT 5054.280 6.800 5057.000 1429.360 ;
    RECT 5059.720 6.800 5062.440 1429.360 ;
    RECT 5065.160 6.800 5067.880 1429.360 ;
    RECT 5070.600 6.800 5073.320 1429.360 ;
    RECT 5076.040 6.800 5078.760 1429.360 ;
    RECT 5081.480 6.800 5084.200 1429.360 ;
    RECT 5086.920 6.800 5089.640 1429.360 ;
    RECT 5092.360 6.800 5095.080 1429.360 ;
    RECT 5097.800 6.800 5100.520 1429.360 ;
    RECT 5103.240 6.800 5105.960 1429.360 ;
    RECT 5108.680 6.800 5111.400 1429.360 ;
    RECT 5114.120 6.800 5116.840 1429.360 ;
    RECT 5119.560 6.800 5122.280 1429.360 ;
    RECT 5125.000 6.800 5127.720 1429.360 ;
    RECT 5130.440 6.800 5133.160 1429.360 ;
    RECT 5135.880 6.800 5138.600 1429.360 ;
    RECT 5141.320 6.800 5144.040 1429.360 ;
    RECT 5146.760 6.800 5149.480 1429.360 ;
    RECT 5152.200 6.800 5154.920 1429.360 ;
    RECT 5157.640 6.800 5160.360 1429.360 ;
    RECT 5163.080 6.800 5165.800 1429.360 ;
    RECT 5168.520 6.800 5171.240 1429.360 ;
    RECT 5173.960 6.800 5176.680 1429.360 ;
    RECT 5179.400 6.800 5182.120 1429.360 ;
    RECT 5184.840 6.800 5187.560 1429.360 ;
    RECT 5190.280 6.800 5193.000 1429.360 ;
    RECT 5195.720 6.800 5198.440 1429.360 ;
    RECT 5201.160 6.800 5203.880 1429.360 ;
    RECT 5206.600 6.800 5209.320 1429.360 ;
    RECT 5212.040 6.800 5214.760 1429.360 ;
    RECT 5217.480 6.800 5220.200 1429.360 ;
    RECT 5222.920 6.800 5225.640 1429.360 ;
    RECT 5228.360 6.800 5231.080 1429.360 ;
    RECT 5233.800 6.800 5236.520 1429.360 ;
    RECT 5239.240 6.800 5241.960 1429.360 ;
    RECT 5244.680 6.800 5247.400 1429.360 ;
    RECT 5250.120 6.800 5252.840 1429.360 ;
    RECT 5255.560 6.800 5258.280 1429.360 ;
    RECT 5261.000 6.800 5263.720 1429.360 ;
    RECT 5266.440 6.800 5269.160 1429.360 ;
    RECT 5271.880 6.800 5274.600 1429.360 ;
    RECT 5277.320 6.800 5280.040 1429.360 ;
    RECT 5282.760 6.800 5285.480 1429.360 ;
    RECT 5288.200 6.800 5290.920 1429.360 ;
    RECT 5293.640 6.800 5296.360 1429.360 ;
    RECT 5299.080 6.800 5301.800 1429.360 ;
    RECT 5304.520 6.800 5307.240 1429.360 ;
    RECT 5309.960 6.800 5312.680 1429.360 ;
    RECT 5315.400 6.800 5318.120 1429.360 ;
    RECT 5320.840 6.800 5323.560 1429.360 ;
    RECT 5326.280 6.800 5329.000 1429.360 ;
    RECT 5331.720 6.800 5334.440 1429.360 ;
    RECT 5337.160 6.800 5339.880 1429.360 ;
    RECT 5342.600 6.800 5345.320 1429.360 ;
    RECT 5348.040 6.800 5350.760 1429.360 ;
    RECT 5353.480 6.800 5356.200 1429.360 ;
    RECT 5358.920 6.800 5361.640 1429.360 ;
    RECT 5364.360 6.800 5367.080 1429.360 ;
    RECT 5369.800 6.800 5372.520 1429.360 ;
    RECT 5375.240 6.800 5377.960 1429.360 ;
    RECT 5380.680 6.800 5383.400 1429.360 ;
    RECT 5386.120 6.800 5388.840 1429.360 ;
    RECT 5391.560 6.800 5394.280 1429.360 ;
    RECT 5397.000 6.800 5399.720 1429.360 ;
    RECT 5402.440 6.800 5405.160 1429.360 ;
    RECT 5407.880 6.800 5410.600 1429.360 ;
    RECT 5413.320 6.800 5416.040 1429.360 ;
    RECT 5418.760 6.800 5421.480 1429.360 ;
    RECT 5424.200 6.800 5426.920 1429.360 ;
    RECT 5429.640 6.800 5432.360 1429.360 ;
    RECT 5435.080 6.800 5437.800 1429.360 ;
    RECT 5440.520 6.800 5443.240 1429.360 ;
    RECT 5445.960 6.800 5448.680 1429.360 ;
    RECT 5451.400 6.800 5454.120 1429.360 ;
    RECT 5456.840 6.800 5459.560 1429.360 ;
    RECT 5462.280 6.800 5465.000 1429.360 ;
    RECT 5467.720 6.800 5470.440 1429.360 ;
    RECT 5473.160 6.800 5475.880 1429.360 ;
    RECT 5478.600 6.800 5481.320 1429.360 ;
    RECT 5484.040 6.800 5486.760 1429.360 ;
    RECT 5489.480 6.800 5492.200 1429.360 ;
    RECT 5494.920 6.800 5497.640 1429.360 ;
    RECT 5500.360 6.800 5503.080 1429.360 ;
    RECT 5505.800 6.800 5508.520 1429.360 ;
    RECT 5511.240 6.800 5513.960 1429.360 ;
    RECT 5516.680 6.800 5519.400 1429.360 ;
    RECT 5522.120 6.800 5524.840 1429.360 ;
    RECT 5527.560 6.800 5530.280 1429.360 ;
    RECT 5533.000 6.800 5535.720 1429.360 ;
    RECT 5538.440 6.800 5541.160 1429.360 ;
    RECT 5543.880 6.800 5546.600 1429.360 ;
    RECT 5549.320 6.800 5552.040 1429.360 ;
    RECT 5554.760 6.800 5557.480 1429.360 ;
    RECT 5560.200 6.800 5562.920 1429.360 ;
    RECT 5565.640 6.800 5568.360 1429.360 ;
    RECT 5571.080 6.800 5573.800 1429.360 ;
    RECT 5576.520 6.800 5579.240 1429.360 ;
    RECT 5581.960 6.800 5584.680 1429.360 ;
    RECT 5587.400 6.800 5590.120 1429.360 ;
    RECT 5592.840 6.800 5595.560 1429.360 ;
    RECT 5598.280 6.800 5601.000 1429.360 ;
    RECT 5603.720 6.800 5606.440 1429.360 ;
    RECT 5609.160 6.800 5611.880 1429.360 ;
    RECT 5614.600 6.800 5617.320 1429.360 ;
    RECT 5620.040 6.800 5622.760 1429.360 ;
    RECT 5625.480 6.800 5628.200 1429.360 ;
    RECT 5630.920 6.800 5633.640 1429.360 ;
    RECT 5636.360 6.800 5639.080 1429.360 ;
    RECT 5641.800 6.800 5644.520 1429.360 ;
    RECT 5647.240 6.800 5649.960 1429.360 ;
    RECT 5652.680 6.800 5655.400 1429.360 ;
    RECT 5658.120 6.800 5660.840 1429.360 ;
    RECT 5663.560 6.800 5666.280 1429.360 ;
    RECT 5669.000 6.800 5671.720 1429.360 ;
    RECT 5674.440 6.800 5677.160 1429.360 ;
    RECT 5679.880 6.800 5682.600 1429.360 ;
    RECT 5685.320 6.800 5688.040 1429.360 ;
    RECT 5690.760 6.800 5693.480 1429.360 ;
    RECT 5696.200 6.800 5698.920 1429.360 ;
    RECT 5701.640 6.800 5704.360 1429.360 ;
    RECT 5707.080 6.800 5709.800 1429.360 ;
    RECT 5712.520 6.800 5715.240 1429.360 ;
    RECT 5717.960 6.800 5720.680 1429.360 ;
    RECT 5723.400 6.800 5726.120 1429.360 ;
    RECT 5728.840 6.800 5731.560 1429.360 ;
    RECT 5734.280 6.800 5737.000 1429.360 ;
    RECT 5739.720 6.800 5742.440 1429.360 ;
    RECT 5745.160 6.800 5747.880 1429.360 ;
    RECT 5750.600 6.800 5753.320 1429.360 ;
    RECT 5756.040 6.800 5758.760 1429.360 ;
    RECT 5761.480 6.800 5764.200 1429.360 ;
    RECT 5766.920 6.800 5769.640 1429.360 ;
    RECT 5772.360 6.800 5775.080 1429.360 ;
    RECT 5777.800 6.800 5780.520 1429.360 ;
    RECT 5783.240 6.800 5785.960 1429.360 ;
    RECT 5788.680 6.800 5791.400 1429.360 ;
    RECT 5794.120 6.800 5796.840 1429.360 ;
    RECT 5799.560 6.800 5802.280 1429.360 ;
    RECT 5805.000 6.800 5807.720 1429.360 ;
    RECT 5810.440 6.800 5813.160 1429.360 ;
    RECT 5815.880 6.800 5818.600 1429.360 ;
    RECT 5821.320 6.800 5824.040 1429.360 ;
    RECT 5826.760 6.800 5829.480 1429.360 ;
    RECT 5832.200 6.800 5834.920 1429.360 ;
    RECT 5837.640 6.800 5840.360 1429.360 ;
    RECT 5843.080 6.800 5845.800 1429.360 ;
    RECT 5848.520 6.800 5851.240 1429.360 ;
    RECT 5853.960 6.800 5856.680 1429.360 ;
    RECT 5859.400 6.800 5862.120 1429.360 ;
    RECT 5864.840 6.800 5871.900 1429.360 ;
    LAYER OVERLAP ;
    RECT 0 0 5871.900 1436.160 ;
  END
END fakeram_512x2048_1r1w

END LIBRARY
