VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_16x52_1r1w
  FOREIGN fakeram_16x52_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 376.280 BY 119.680 ;
  CLASS BLOCK ;
  PIN w0_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 6.650 0.800 6.950 ;
    END
  END w0_mask_in[0]
  PIN w0_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 9.370 0.800 9.670 ;
    END
  END w0_mask_in[1]
  PIN w0_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 12.090 0.800 12.390 ;
    END
  END w0_mask_in[2]
  PIN w0_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.810 0.800 15.110 ;
    END
  END w0_mask_in[3]
  PIN w0_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 17.530 0.800 17.830 ;
    END
  END w0_mask_in[4]
  PIN w0_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.250 0.800 20.550 ;
    END
  END w0_mask_in[5]
  PIN w0_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.970 0.800 23.270 ;
    END
  END w0_mask_in[6]
  PIN w0_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 25.690 0.800 25.990 ;
    END
  END w0_mask_in[7]
  PIN w0_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 28.410 0.800 28.710 ;
    END
  END w0_mask_in[8]
  PIN w0_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.130 0.800 31.430 ;
    END
  END w0_mask_in[9]
  PIN w0_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 33.850 0.800 34.150 ;
    END
  END w0_mask_in[10]
  PIN w0_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 36.570 0.800 36.870 ;
    END
  END w0_mask_in[11]
  PIN w0_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.290 0.800 39.590 ;
    END
  END w0_mask_in[12]
  PIN w0_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 42.010 0.800 42.310 ;
    END
  END w0_mask_in[13]
  PIN w0_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 44.730 0.800 45.030 ;
    END
  END w0_mask_in[14]
  PIN w0_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 47.450 0.800 47.750 ;
    END
  END w0_mask_in[15]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 56.970 0.800 57.270 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 59.690 0.800 59.990 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 62.410 0.800 62.710 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 65.130 0.800 65.430 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.850 0.800 68.150 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 70.570 0.800 70.870 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 73.290 0.800 73.590 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.010 0.800 76.310 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 78.730 0.800 79.030 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 81.450 0.800 81.750 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 84.170 0.800 84.470 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 86.890 0.800 87.190 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.610 0.800 89.910 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 92.330 0.800 92.630 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 95.050 0.800 95.350 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 97.770 0.800 98.070 ;
    END
  END w0_wd_in[15]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 0.000 4.670 0.350 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 27.070 0.000 27.210 0.350 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 49.610 0.000 49.750 0.350 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 72.150 0.000 72.290 0.350 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 94.690 0.000 94.830 0.350 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 117.230 0.000 117.370 0.350 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 139.770 0.000 139.910 0.350 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 162.310 0.000 162.450 0.350 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 184.850 0.000 184.990 0.350 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 207.390 0.000 207.530 0.350 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 229.930 0.000 230.070 0.350 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 252.470 0.000 252.610 0.350 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 275.010 0.000 275.150 0.350 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 297.550 0.000 297.690 0.350 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 320.090 0.000 320.230 0.350 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 342.630 0.000 342.770 0.350 ;
    END
  END r0_rd_out[15]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 6.650 376.280 6.950 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 12.090 376.280 12.390 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 17.530 376.280 17.830 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 22.970 376.280 23.270 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 28.410 376.280 28.710 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 33.850 376.280 34.150 ;
    END
  END w0_addr_in[5]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 119.330 4.670 119.680 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 24.770 119.330 24.910 119.680 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 45.010 119.330 45.150 119.680 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 65.250 119.330 65.390 119.680 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 85.490 119.330 85.630 119.680 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 105.730 119.330 105.870 119.680 ;
    END
  END r0_addr_in[5]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 35.210 376.280 35.510 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 36.570 376.280 36.870 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 37.930 376.280 38.230 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 106.650 119.330 106.790 119.680 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 107.570 119.330 107.710 119.680 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 3.240 6.800 5.960 112.880 ;
      RECT 14.120 6.800 16.840 112.880 ;
      RECT 25.000 6.800 27.720 112.880 ;
      RECT 35.880 6.800 38.600 112.880 ;
      RECT 46.760 6.800 49.480 112.880 ;
      RECT 57.640 6.800 60.360 112.880 ;
      RECT 68.520 6.800 71.240 112.880 ;
      RECT 79.400 6.800 82.120 112.880 ;
      RECT 90.280 6.800 93.000 112.880 ;
      RECT 101.160 6.800 103.880 112.880 ;
      RECT 112.040 6.800 114.760 112.880 ;
      RECT 122.920 6.800 125.640 112.880 ;
      RECT 133.800 6.800 136.520 112.880 ;
      RECT 144.680 6.800 147.400 112.880 ;
      RECT 155.560 6.800 158.280 112.880 ;
      RECT 166.440 6.800 169.160 112.880 ;
      RECT 177.320 6.800 180.040 112.880 ;
      RECT 188.200 6.800 190.920 112.880 ;
      RECT 199.080 6.800 201.800 112.880 ;
      RECT 209.960 6.800 212.680 112.880 ;
      RECT 220.840 6.800 223.560 112.880 ;
      RECT 231.720 6.800 234.440 112.880 ;
      RECT 242.600 6.800 245.320 112.880 ;
      RECT 253.480 6.800 256.200 112.880 ;
      RECT 264.360 6.800 267.080 112.880 ;
      RECT 275.240 6.800 277.960 112.880 ;
      RECT 286.120 6.800 288.840 112.880 ;
      RECT 297.000 6.800 299.720 112.880 ;
      RECT 307.880 6.800 310.600 112.880 ;
      RECT 318.760 6.800 321.480 112.880 ;
      RECT 329.640 6.800 332.360 112.880 ;
      RECT 340.520 6.800 343.240 112.880 ;
      RECT 351.400 6.800 354.120 112.880 ;
      RECT 362.280 6.800 365.000 112.880 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 8.680 6.800 11.400 112.880 ;
      RECT 19.560 6.800 22.280 112.880 ;
      RECT 30.440 6.800 33.160 112.880 ;
      RECT 41.320 6.800 44.040 112.880 ;
      RECT 52.200 6.800 54.920 112.880 ;
      RECT 63.080 6.800 65.800 112.880 ;
      RECT 73.960 6.800 76.680 112.880 ;
      RECT 84.840 6.800 87.560 112.880 ;
      RECT 95.720 6.800 98.440 112.880 ;
      RECT 106.600 6.800 109.320 112.880 ;
      RECT 117.480 6.800 120.200 112.880 ;
      RECT 128.360 6.800 131.080 112.880 ;
      RECT 139.240 6.800 141.960 112.880 ;
      RECT 150.120 6.800 152.840 112.880 ;
      RECT 161.000 6.800 163.720 112.880 ;
      RECT 171.880 6.800 174.600 112.880 ;
      RECT 182.760 6.800 185.480 112.880 ;
      RECT 193.640 6.800 196.360 112.880 ;
      RECT 204.520 6.800 207.240 112.880 ;
      RECT 215.400 6.800 218.120 112.880 ;
      RECT 226.280 6.800 229.000 112.880 ;
      RECT 237.160 6.800 239.880 112.880 ;
      RECT 248.040 6.800 250.760 112.880 ;
      RECT 258.920 6.800 261.640 112.880 ;
      RECT 269.800 6.800 272.520 112.880 ;
      RECT 280.680 6.800 283.400 112.880 ;
      RECT 291.560 6.800 294.280 112.880 ;
      RECT 302.440 6.800 305.160 112.880 ;
      RECT 313.320 6.800 316.040 112.880 ;
      RECT 324.200 6.800 326.920 112.880 ;
      RECT 335.080 6.800 337.800 112.880 ;
      RECT 345.960 6.800 348.680 112.880 ;
      RECT 356.840 6.800 359.560 112.880 ;
      RECT 367.720 6.800 370.440 112.880 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 376.280 119.680 ;
    LAYER met2 ;
    RECT 0 0 376.280 119.680 ;
    LAYER met3 ;
    RECT 0.800 0 376.280 119.680 ;
    LAYER met4 ;
    RECT 0 0 376.280 6.800 ;
    RECT 0 112.880 376.280 119.680 ;
    RECT 0.000 6.800 3.240 112.880 ;
    RECT 5.960 6.800 8.680 112.880 ;
    RECT 11.400 6.800 14.120 112.880 ;
    RECT 16.840 6.800 19.560 112.880 ;
    RECT 22.280 6.800 25.000 112.880 ;
    RECT 27.720 6.800 30.440 112.880 ;
    RECT 33.160 6.800 35.880 112.880 ;
    RECT 38.600 6.800 41.320 112.880 ;
    RECT 44.040 6.800 46.760 112.880 ;
    RECT 49.480 6.800 52.200 112.880 ;
    RECT 54.920 6.800 57.640 112.880 ;
    RECT 60.360 6.800 63.080 112.880 ;
    RECT 65.800 6.800 68.520 112.880 ;
    RECT 71.240 6.800 73.960 112.880 ;
    RECT 76.680 6.800 79.400 112.880 ;
    RECT 82.120 6.800 84.840 112.880 ;
    RECT 87.560 6.800 90.280 112.880 ;
    RECT 93.000 6.800 95.720 112.880 ;
    RECT 98.440 6.800 101.160 112.880 ;
    RECT 103.880 6.800 106.600 112.880 ;
    RECT 109.320 6.800 112.040 112.880 ;
    RECT 114.760 6.800 117.480 112.880 ;
    RECT 120.200 6.800 122.920 112.880 ;
    RECT 125.640 6.800 128.360 112.880 ;
    RECT 131.080 6.800 133.800 112.880 ;
    RECT 136.520 6.800 139.240 112.880 ;
    RECT 141.960 6.800 144.680 112.880 ;
    RECT 147.400 6.800 150.120 112.880 ;
    RECT 152.840 6.800 155.560 112.880 ;
    RECT 158.280 6.800 161.000 112.880 ;
    RECT 163.720 6.800 166.440 112.880 ;
    RECT 169.160 6.800 171.880 112.880 ;
    RECT 174.600 6.800 177.320 112.880 ;
    RECT 180.040 6.800 182.760 112.880 ;
    RECT 185.480 6.800 188.200 112.880 ;
    RECT 190.920 6.800 193.640 112.880 ;
    RECT 196.360 6.800 199.080 112.880 ;
    RECT 201.800 6.800 204.520 112.880 ;
    RECT 207.240 6.800 209.960 112.880 ;
    RECT 212.680 6.800 215.400 112.880 ;
    RECT 218.120 6.800 220.840 112.880 ;
    RECT 223.560 6.800 226.280 112.880 ;
    RECT 229.000 6.800 231.720 112.880 ;
    RECT 234.440 6.800 237.160 112.880 ;
    RECT 239.880 6.800 242.600 112.880 ;
    RECT 245.320 6.800 248.040 112.880 ;
    RECT 250.760 6.800 253.480 112.880 ;
    RECT 256.200 6.800 258.920 112.880 ;
    RECT 261.640 6.800 264.360 112.880 ;
    RECT 267.080 6.800 269.800 112.880 ;
    RECT 272.520 6.800 275.240 112.880 ;
    RECT 277.960 6.800 280.680 112.880 ;
    RECT 283.400 6.800 286.120 112.880 ;
    RECT 288.840 6.800 291.560 112.880 ;
    RECT 294.280 6.800 297.000 112.880 ;
    RECT 299.720 6.800 302.440 112.880 ;
    RECT 305.160 6.800 307.880 112.880 ;
    RECT 310.600 6.800 313.320 112.880 ;
    RECT 316.040 6.800 318.760 112.880 ;
    RECT 321.480 6.800 324.200 112.880 ;
    RECT 326.920 6.800 329.640 112.880 ;
    RECT 332.360 6.800 335.080 112.880 ;
    RECT 337.800 6.800 340.520 112.880 ;
    RECT 343.240 6.800 345.960 112.880 ;
    RECT 348.680 6.800 351.400 112.880 ;
    RECT 354.120 6.800 356.840 112.880 ;
    RECT 359.560 6.800 362.280 112.880 ;
    RECT 365.000 6.800 367.720 112.880 ;
    RECT 370.440 6.800 376.280 112.880 ;
    LAYER OVERLAP ;
    RECT 0 0 376.280 119.680 ;
  END
END fakeram_16x52_1r1w

END LIBRARY
