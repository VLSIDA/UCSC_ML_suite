VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_512x2048_1r1w
  FOREIGN fakeram_512x2048_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 78.660 BY 229.600 ;
  CLASS BLOCK ;
  PIN w_mask_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 -0.035 0.070 0.035 ;
    END
  END w_mask_w1[0]
  PIN w_mask_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_w1[1]
  PIN w_mask_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_w1[2]
  PIN w_mask_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_w1[3]
  PIN w_mask_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_w1[4]
  PIN w_mask_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_w1[5]
  PIN w_mask_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_w1[6]
  PIN w_mask_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END w_mask_w1[7]
  PIN w_mask_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_w1[8]
  PIN w_mask_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END w_mask_w1[9]
  PIN w_mask_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END w_mask_w1[10]
  PIN w_mask_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END w_mask_w1[11]
  PIN w_mask_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END w_mask_w1[12]
  PIN w_mask_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END w_mask_w1[13]
  PIN w_mask_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END w_mask_w1[14]
  PIN w_mask_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END w_mask_w1[15]
  PIN w_mask_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END w_mask_w1[16]
  PIN w_mask_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END w_mask_w1[17]
  PIN rd_out_r1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.045 0.070 59.115 ;
    END
  END rd_out_r1[0]
  PIN rd_out_r1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.405 0.070 62.475 ;
    END
  END rd_out_r1[1]
  PIN rd_out_r1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.765 0.070 65.835 ;
    END
  END rd_out_r1[2]
  PIN rd_out_r1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.125 0.070 69.195 ;
    END
  END rd_out_r1[3]
  PIN rd_out_r1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.485 0.070 72.555 ;
    END
  END rd_out_r1[4]
  PIN rd_out_r1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.845 0.070 75.915 ;
    END
  END rd_out_r1[5]
  PIN rd_out_r1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.205 0.070 79.275 ;
    END
  END rd_out_r1[6]
  PIN rd_out_r1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.565 0.070 82.635 ;
    END
  END rd_out_r1[7]
  PIN rd_out_r1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.925 0.070 85.995 ;
    END
  END rd_out_r1[8]
  PIN rd_out_r1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.285 0.070 89.355 ;
    END
  END rd_out_r1[9]
  PIN rd_out_r1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.645 0.070 92.715 ;
    END
  END rd_out_r1[10]
  PIN rd_out_r1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.005 0.070 96.075 ;
    END
  END rd_out_r1[11]
  PIN rd_out_r1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.365 0.070 99.435 ;
    END
  END rd_out_r1[12]
  PIN rd_out_r1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.725 0.070 102.795 ;
    END
  END rd_out_r1[13]
  PIN rd_out_r1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.085 0.070 106.155 ;
    END
  END rd_out_r1[14]
  PIN rd_out_r1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.445 0.070 109.515 ;
    END
  END rd_out_r1[15]
  PIN rd_out_r1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.805 0.070 112.875 ;
    END
  END rd_out_r1[16]
  PIN rd_out_r1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.165 0.070 116.235 ;
    END
  END rd_out_r1[17]
  PIN wd_in_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.125 0.070 118.195 ;
    END
  END wd_in_w1[0]
  PIN wd_in_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.485 0.070 121.555 ;
    END
  END wd_in_w1[1]
  PIN wd_in_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.845 0.070 124.915 ;
    END
  END wd_in_w1[2]
  PIN wd_in_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.205 0.070 128.275 ;
    END
  END wd_in_w1[3]
  PIN wd_in_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.565 0.070 131.635 ;
    END
  END wd_in_w1[4]
  PIN wd_in_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.925 0.070 134.995 ;
    END
  END wd_in_w1[5]
  PIN wd_in_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.285 0.070 138.355 ;
    END
  END wd_in_w1[6]
  PIN wd_in_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.645 0.070 141.715 ;
    END
  END wd_in_w1[7]
  PIN wd_in_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.005 0.070 145.075 ;
    END
  END wd_in_w1[8]
  PIN wd_in_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.365 0.070 148.435 ;
    END
  END wd_in_w1[9]
  PIN wd_in_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.725 0.070 151.795 ;
    END
  END wd_in_w1[10]
  PIN wd_in_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.085 0.070 155.155 ;
    END
  END wd_in_w1[11]
  PIN wd_in_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.445 0.070 158.515 ;
    END
  END wd_in_w1[12]
  PIN wd_in_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.805 0.070 161.875 ;
    END
  END wd_in_w1[13]
  PIN wd_in_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.165 0.070 165.235 ;
    END
  END wd_in_w1[14]
  PIN wd_in_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.525 0.070 168.595 ;
    END
  END wd_in_w1[15]
  PIN wd_in_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.885 0.070 171.955 ;
    END
  END wd_in_w1[16]
  PIN wd_in_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.245 0.070 175.315 ;
    END
  END wd_in_w1[17]
  PIN addr_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.205 0.070 177.275 ;
    END
  END addr_w1[0]
  PIN addr_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.565 0.070 180.635 ;
    END
  END addr_w1[1]
  PIN addr_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.925 0.070 183.995 ;
    END
  END addr_w1[2]
  PIN addr_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.285 0.070 187.355 ;
    END
  END addr_w1[3]
  PIN addr_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.645 0.070 190.715 ;
    END
  END addr_w1[4]
  PIN addr_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.005 0.070 194.075 ;
    END
  END addr_w1[5]
  PIN addr_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.365 0.070 197.435 ;
    END
  END addr_w1[6]
  PIN addr_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.725 0.070 200.795 ;
    END
  END addr_w1[7]
  PIN addr_r1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.685 0.070 202.755 ;
    END
  END addr_r1[0]
  PIN addr_r1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.045 0.070 206.115 ;
    END
  END addr_r1[1]
  PIN addr_r1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.405 0.070 209.475 ;
    END
  END addr_r1[2]
  PIN addr_r1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.765 0.070 212.835 ;
    END
  END addr_r1[3]
  PIN addr_r1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.125 0.070 216.195 ;
    END
  END addr_r1[4]
  PIN addr_r1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.485 0.070 219.555 ;
    END
  END addr_r1[5]
  PIN addr_r1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.845 0.070 222.915 ;
    END
  END addr_r1[6]
  PIN addr_r1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.205 0.070 226.275 ;
    END
  END addr_r1[7]
  PIN we_in_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.165 0.070 228.235 ;
    END
  END we_in_w1
  PIN ce_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.725 0.070 228.795 ;
    END
  END ce_w1
  PIN ce_r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.685 0.070 230.755 ;
    END
  END ce_r1
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.645 0.070 232.715 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 228.200 ;
      RECT 3.500 1.400 3.780 228.200 ;
      RECT 5.740 1.400 6.020 228.200 ;
      RECT 7.980 1.400 8.260 228.200 ;
      RECT 10.220 1.400 10.500 228.200 ;
      RECT 12.460 1.400 12.740 228.200 ;
      RECT 14.700 1.400 14.980 228.200 ;
      RECT 16.940 1.400 17.220 228.200 ;
      RECT 19.180 1.400 19.460 228.200 ;
      RECT 21.420 1.400 21.700 228.200 ;
      RECT 23.660 1.400 23.940 228.200 ;
      RECT 25.900 1.400 26.180 228.200 ;
      RECT 28.140 1.400 28.420 228.200 ;
      RECT 30.380 1.400 30.660 228.200 ;
      RECT 32.620 1.400 32.900 228.200 ;
      RECT 34.860 1.400 35.140 228.200 ;
      RECT 37.100 1.400 37.380 228.200 ;
      RECT 39.340 1.400 39.620 228.200 ;
      RECT 41.580 1.400 41.860 228.200 ;
      RECT 43.820 1.400 44.100 228.200 ;
      RECT 46.060 1.400 46.340 228.200 ;
      RECT 48.300 1.400 48.580 228.200 ;
      RECT 50.540 1.400 50.820 228.200 ;
      RECT 52.780 1.400 53.060 228.200 ;
      RECT 55.020 1.400 55.300 228.200 ;
      RECT 57.260 1.400 57.540 228.200 ;
      RECT 59.500 1.400 59.780 228.200 ;
      RECT 61.740 1.400 62.020 228.200 ;
      RECT 63.980 1.400 64.260 228.200 ;
      RECT 66.220 1.400 66.500 228.200 ;
      RECT 68.460 1.400 68.740 228.200 ;
      RECT 70.700 1.400 70.980 228.200 ;
      RECT 72.940 1.400 73.220 228.200 ;
      RECT 75.180 1.400 75.460 228.200 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 228.200 ;
      RECT 4.620 1.400 4.900 228.200 ;
      RECT 6.860 1.400 7.140 228.200 ;
      RECT 9.100 1.400 9.380 228.200 ;
      RECT 11.340 1.400 11.620 228.200 ;
      RECT 13.580 1.400 13.860 228.200 ;
      RECT 15.820 1.400 16.100 228.200 ;
      RECT 18.060 1.400 18.340 228.200 ;
      RECT 20.300 1.400 20.580 228.200 ;
      RECT 22.540 1.400 22.820 228.200 ;
      RECT 24.780 1.400 25.060 228.200 ;
      RECT 27.020 1.400 27.300 228.200 ;
      RECT 29.260 1.400 29.540 228.200 ;
      RECT 31.500 1.400 31.780 228.200 ;
      RECT 33.740 1.400 34.020 228.200 ;
      RECT 35.980 1.400 36.260 228.200 ;
      RECT 38.220 1.400 38.500 228.200 ;
      RECT 40.460 1.400 40.740 228.200 ;
      RECT 42.700 1.400 42.980 228.200 ;
      RECT 44.940 1.400 45.220 228.200 ;
      RECT 47.180 1.400 47.460 228.200 ;
      RECT 49.420 1.400 49.700 228.200 ;
      RECT 51.660 1.400 51.940 228.200 ;
      RECT 53.900 1.400 54.180 228.200 ;
      RECT 56.140 1.400 56.420 228.200 ;
      RECT 58.380 1.400 58.660 228.200 ;
      RECT 60.620 1.400 60.900 228.200 ;
      RECT 62.860 1.400 63.140 228.200 ;
      RECT 65.100 1.400 65.380 228.200 ;
      RECT 67.340 1.400 67.620 228.200 ;
      RECT 69.580 1.400 69.860 228.200 ;
      RECT 71.820 1.400 72.100 228.200 ;
      RECT 74.060 1.400 74.340 228.200 ;
      RECT 76.300 1.400 76.580 228.200 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 78.660 229.600 ;
    LAYER metal2 ;
    RECT 0 0 78.660 229.600 ;
    LAYER metal3 ;
    RECT 0.070 0 78.660 229.600 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 4.725 ;
    RECT 0 4.795 0.070 8.085 ;
    RECT 0 8.155 0.070 11.445 ;
    RECT 0 11.515 0.070 14.805 ;
    RECT 0 14.875 0.070 18.165 ;
    RECT 0 18.235 0.070 21.525 ;
    RECT 0 21.595 0.070 24.885 ;
    RECT 0 24.955 0.070 28.245 ;
    RECT 0 28.315 0.070 31.605 ;
    RECT 0 31.675 0.070 34.965 ;
    RECT 0 35.035 0.070 38.325 ;
    RECT 0 38.395 0.070 41.685 ;
    RECT 0 41.755 0.070 45.045 ;
    RECT 0 45.115 0.070 48.405 ;
    RECT 0 48.475 0.070 51.765 ;
    RECT 0 51.835 0.070 55.125 ;
    RECT 0 55.195 0.070 58.485 ;
    RECT 0 58.555 0.070 60.445 ;
    RECT 0 60.515 0.070 63.805 ;
    RECT 0 63.875 0.070 67.165 ;
    RECT 0 67.235 0.070 70.525 ;
    RECT 0 70.595 0.070 73.885 ;
    RECT 0 73.955 0.070 77.245 ;
    RECT 0 77.315 0.070 80.605 ;
    RECT 0 80.675 0.070 83.965 ;
    RECT 0 84.035 0.070 87.325 ;
    RECT 0 87.395 0.070 90.685 ;
    RECT 0 90.755 0.070 94.045 ;
    RECT 0 94.115 0.070 97.405 ;
    RECT 0 97.475 0.070 100.765 ;
    RECT 0 100.835 0.070 104.125 ;
    RECT 0 104.195 0.070 107.485 ;
    RECT 0 107.555 0.070 110.845 ;
    RECT 0 110.915 0.070 114.205 ;
    RECT 0 114.275 0.070 117.565 ;
    RECT 0 117.635 0.070 119.525 ;
    RECT 0 119.595 0.070 122.885 ;
    RECT 0 122.955 0.070 126.245 ;
    RECT 0 126.315 0.070 129.605 ;
    RECT 0 129.675 0.070 132.965 ;
    RECT 0 133.035 0.070 136.325 ;
    RECT 0 136.395 0.070 139.685 ;
    RECT 0 139.755 0.070 143.045 ;
    RECT 0 143.115 0.070 146.405 ;
    RECT 0 146.475 0.070 149.765 ;
    RECT 0 149.835 0.070 153.125 ;
    RECT 0 153.195 0.070 156.485 ;
    RECT 0 156.555 0.070 159.845 ;
    RECT 0 159.915 0.070 163.205 ;
    RECT 0 163.275 0.070 166.565 ;
    RECT 0 166.635 0.070 169.925 ;
    RECT 0 169.995 0.070 173.285 ;
    RECT 0 173.355 0.070 176.645 ;
    RECT 0 176.715 0.070 178.605 ;
    RECT 0 178.675 0.070 181.965 ;
    RECT 0 182.035 0.070 185.325 ;
    RECT 0 185.395 0.070 188.685 ;
    RECT 0 188.755 0.070 192.045 ;
    RECT 0 192.115 0.070 195.405 ;
    RECT 0 195.475 0.070 198.765 ;
    RECT 0 198.835 0.070 202.125 ;
    RECT 0 202.195 0.070 204.085 ;
    RECT 0 204.155 0.070 207.445 ;
    RECT 0 207.515 0.070 210.805 ;
    RECT 0 210.875 0.070 229.600 ;
    LAYER metal4 ;
    RECT 0 0 78.660 1.400 ;
    RECT 0 228.200 78.660 229.600 ;
    RECT 0.000 1.400 1.260 228.200 ;
    RECT 1.540 1.400 2.380 228.200 ;
    RECT 2.660 1.400 3.500 228.200 ;
    RECT 3.780 1.400 4.620 228.200 ;
    RECT 4.900 1.400 5.740 228.200 ;
    RECT 6.020 1.400 6.860 228.200 ;
    RECT 7.140 1.400 7.980 228.200 ;
    RECT 8.260 1.400 9.100 228.200 ;
    RECT 9.380 1.400 10.220 228.200 ;
    RECT 10.500 1.400 11.340 228.200 ;
    RECT 11.620 1.400 12.460 228.200 ;
    RECT 12.740 1.400 13.580 228.200 ;
    RECT 13.860 1.400 14.700 228.200 ;
    RECT 14.980 1.400 15.820 228.200 ;
    RECT 16.100 1.400 16.940 228.200 ;
    RECT 17.220 1.400 18.060 228.200 ;
    RECT 18.340 1.400 19.180 228.200 ;
    RECT 19.460 1.400 20.300 228.200 ;
    RECT 20.580 1.400 21.420 228.200 ;
    RECT 21.700 1.400 22.540 228.200 ;
    RECT 22.820 1.400 23.660 228.200 ;
    RECT 23.940 1.400 24.780 228.200 ;
    RECT 25.060 1.400 25.900 228.200 ;
    RECT 26.180 1.400 27.020 228.200 ;
    RECT 27.300 1.400 28.140 228.200 ;
    RECT 28.420 1.400 29.260 228.200 ;
    RECT 29.540 1.400 30.380 228.200 ;
    RECT 30.660 1.400 31.500 228.200 ;
    RECT 31.780 1.400 32.620 228.200 ;
    RECT 32.900 1.400 33.740 228.200 ;
    RECT 34.020 1.400 34.860 228.200 ;
    RECT 35.140 1.400 35.980 228.200 ;
    RECT 36.260 1.400 37.100 228.200 ;
    RECT 37.380 1.400 38.220 228.200 ;
    RECT 38.500 1.400 39.340 228.200 ;
    RECT 39.620 1.400 40.460 228.200 ;
    RECT 40.740 1.400 41.580 228.200 ;
    RECT 41.860 1.400 42.700 228.200 ;
    RECT 42.980 1.400 43.820 228.200 ;
    RECT 44.100 1.400 44.940 228.200 ;
    RECT 45.220 1.400 46.060 228.200 ;
    RECT 46.340 1.400 47.180 228.200 ;
    RECT 47.460 1.400 48.300 228.200 ;
    RECT 48.580 1.400 49.420 228.200 ;
    RECT 49.700 1.400 50.540 228.200 ;
    RECT 50.820 1.400 51.660 228.200 ;
    RECT 51.940 1.400 52.780 228.200 ;
    RECT 53.060 1.400 53.900 228.200 ;
    RECT 54.180 1.400 55.020 228.200 ;
    RECT 55.300 1.400 56.140 228.200 ;
    RECT 56.420 1.400 57.260 228.200 ;
    RECT 57.540 1.400 58.380 228.200 ;
    RECT 58.660 1.400 59.500 228.200 ;
    RECT 59.780 1.400 60.620 228.200 ;
    RECT 60.900 1.400 61.740 228.200 ;
    RECT 62.020 1.400 62.860 228.200 ;
    RECT 63.140 1.400 63.980 228.200 ;
    RECT 64.260 1.400 65.100 228.200 ;
    RECT 65.380 1.400 66.220 228.200 ;
    RECT 66.500 1.400 67.340 228.200 ;
    RECT 67.620 1.400 68.460 228.200 ;
    RECT 68.740 1.400 69.580 228.200 ;
    RECT 69.860 1.400 70.700 228.200 ;
    RECT 70.980 1.400 71.820 228.200 ;
    RECT 72.100 1.400 72.940 228.200 ;
    RECT 73.220 1.400 74.060 228.200 ;
    RECT 74.340 1.400 75.180 228.200 ;
    RECT 75.460 1.400 76.300 228.200 ;
    RECT 76.580 1.400 78.660 228.200 ;
    LAYER OVERLAP ;
    RECT 0 0 78.660 229.600 ;
  END
END fakeram_512x2048_1r1w

END LIBRARY
