VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_20x64_2r1w
  FOREIGN fakeram_20x64_2r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 98.990 BY 134.400 ;
  CLASS BLOCK ;
  PIN w_mask_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 0.945 0.070 1.015 ;
    END
  END w_mask_w1[0]
  PIN w_mask_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_w1[1]
  PIN w_mask_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_w1[2]
  PIN w_mask_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_w1[3]
  PIN w_mask_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.225 0.070 8.295 ;
    END
  END w_mask_w1[4]
  PIN w_mask_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_w1[5]
  PIN w_mask_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.865 0.070 11.935 ;
    END
  END w_mask_w1[6]
  PIN w_mask_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.685 0.070 13.755 ;
    END
  END w_mask_w1[7]
  PIN w_mask_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_w1[8]
  PIN w_mask_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.325 0.070 17.395 ;
    END
  END w_mask_w1[9]
  PIN w_mask_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.145 0.070 19.215 ;
    END
  END w_mask_w1[10]
  PIN w_mask_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_w1[11]
  PIN w_mask_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.785 0.070 22.855 ;
    END
  END w_mask_w1[12]
  PIN w_mask_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.605 0.070 24.675 ;
    END
  END w_mask_w1[13]
  PIN w_mask_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END w_mask_w1[14]
  PIN w_mask_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.245 0.070 28.315 ;
    END
  END w_mask_w1[15]
  PIN w_mask_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.065 0.070 30.135 ;
    END
  END w_mask_w1[16]
  PIN w_mask_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END w_mask_w1[17]
  PIN w_mask_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.705 0.070 33.775 ;
    END
  END w_mask_w1[18]
  PIN w_mask_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.525 0.070 35.595 ;
    END
  END w_mask_w1[19]
  PIN rd_out_r1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END rd_out_r1[0]
  PIN rd_out_r1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.745 0.070 38.815 ;
    END
  END rd_out_r1[1]
  PIN rd_out_r1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END rd_out_r1[2]
  PIN rd_out_r1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END rd_out_r1[3]
  PIN rd_out_r1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.205 0.070 44.275 ;
    END
  END rd_out_r1[4]
  PIN rd_out_r1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.025 0.070 46.095 ;
    END
  END rd_out_r1[5]
  PIN rd_out_r1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out_r1[6]
  PIN rd_out_r1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.665 0.070 49.735 ;
    END
  END rd_out_r1[7]
  PIN rd_out_r1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.485 0.070 51.555 ;
    END
  END rd_out_r1[8]
  PIN rd_out_r1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END rd_out_r1[9]
  PIN rd_out_r1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.125 0.070 55.195 ;
    END
  END rd_out_r1[10]
  PIN rd_out_r1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.945 0.070 57.015 ;
    END
  END rd_out_r1[11]
  PIN rd_out_r1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END rd_out_r1[12]
  PIN rd_out_r1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.585 0.070 60.655 ;
    END
  END rd_out_r1[13]
  PIN rd_out_r1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.405 0.070 62.475 ;
    END
  END rd_out_r1[14]
  PIN rd_out_r1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END rd_out_r1[15]
  PIN rd_out_r1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.045 0.070 66.115 ;
    END
  END rd_out_r1[16]
  PIN rd_out_r1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.865 0.070 67.935 ;
    END
  END rd_out_r1[17]
  PIN rd_out_r1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END rd_out_r1[18]
  PIN rd_out_r1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.505 0.070 71.575 ;
    END
  END rd_out_r1[19]
  PIN rd_out_r2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.905 0.070 72.975 ;
    END
  END rd_out_r2[0]
  PIN rd_out_r2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END rd_out_r2[1]
  PIN rd_out_r2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.545 0.070 76.615 ;
    END
  END rd_out_r2[2]
  PIN rd_out_r2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.365 0.070 78.435 ;
    END
  END rd_out_r2[3]
  PIN rd_out_r2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END rd_out_r2[4]
  PIN rd_out_r2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.005 0.070 82.075 ;
    END
  END rd_out_r2[5]
  PIN rd_out_r2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.825 0.070 83.895 ;
    END
  END rd_out_r2[6]
  PIN rd_out_r2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END rd_out_r2[7]
  PIN rd_out_r2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.465 0.070 87.535 ;
    END
  END rd_out_r2[8]
  PIN rd_out_r2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.285 0.070 89.355 ;
    END
  END rd_out_r2[9]
  PIN rd_out_r2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.105 0.070 91.175 ;
    END
  END rd_out_r2[10]
  PIN rd_out_r2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.925 0.070 92.995 ;
    END
  END rd_out_r2[11]
  PIN rd_out_r2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.745 0.070 94.815 ;
    END
  END rd_out_r2[12]
  PIN rd_out_r2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.565 0.070 96.635 ;
    END
  END rd_out_r2[13]
  PIN rd_out_r2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.385 0.070 98.455 ;
    END
  END rd_out_r2[14]
  PIN rd_out_r2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.205 0.070 100.275 ;
    END
  END rd_out_r2[15]
  PIN rd_out_r2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.025 0.070 102.095 ;
    END
  END rd_out_r2[16]
  PIN rd_out_r2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.845 0.070 103.915 ;
    END
  END rd_out_r2[17]
  PIN rd_out_r2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.665 0.070 105.735 ;
    END
  END rd_out_r2[18]
  PIN rd_out_r2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.485 0.070 107.555 ;
    END
  END rd_out_r2[19]
  PIN wd_in_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.885 0.070 108.955 ;
    END
  END wd_in_w1[0]
  PIN wd_in_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.705 0.070 110.775 ;
    END
  END wd_in_w1[1]
  PIN wd_in_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.525 0.070 112.595 ;
    END
  END wd_in_w1[2]
  PIN wd_in_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.345 0.070 114.415 ;
    END
  END wd_in_w1[3]
  PIN wd_in_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.165 0.070 116.235 ;
    END
  END wd_in_w1[4]
  PIN wd_in_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.985 0.070 118.055 ;
    END
  END wd_in_w1[5]
  PIN wd_in_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.805 0.070 119.875 ;
    END
  END wd_in_w1[6]
  PIN wd_in_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.625 0.070 121.695 ;
    END
  END wd_in_w1[7]
  PIN wd_in_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.445 0.070 123.515 ;
    END
  END wd_in_w1[8]
  PIN wd_in_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.265 0.070 125.335 ;
    END
  END wd_in_w1[9]
  PIN wd_in_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.085 0.070 127.155 ;
    END
  END wd_in_w1[10]
  PIN wd_in_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.905 0.070 128.975 ;
    END
  END wd_in_w1[11]
  PIN wd_in_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.725 0.070 130.795 ;
    END
  END wd_in_w1[12]
  PIN wd_in_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.545 0.070 132.615 ;
    END
  END wd_in_w1[13]
  PIN wd_in_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.365 0.070 134.435 ;
    END
  END wd_in_w1[14]
  PIN wd_in_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.185 0.070 136.255 ;
    END
  END wd_in_w1[15]
  PIN wd_in_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.005 0.070 138.075 ;
    END
  END wd_in_w1[16]
  PIN wd_in_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.825 0.070 139.895 ;
    END
  END wd_in_w1[17]
  PIN wd_in_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.645 0.070 141.715 ;
    END
  END wd_in_w1[18]
  PIN wd_in_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.465 0.070 143.535 ;
    END
  END wd_in_w1[19]
  PIN addr_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.865 0.070 144.935 ;
    END
  END addr_w1[0]
  PIN addr_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.685 0.070 146.755 ;
    END
  END addr_w1[1]
  PIN addr_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.505 0.070 148.575 ;
    END
  END addr_w1[2]
  PIN addr_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.325 0.070 150.395 ;
    END
  END addr_w1[3]
  PIN addr_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.145 0.070 152.215 ;
    END
  END addr_w1[4]
  PIN addr_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.965 0.070 154.035 ;
    END
  END addr_w1[5]
  PIN addr_r1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.365 0.070 155.435 ;
    END
  END addr_r1[0]
  PIN addr_r1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.185 0.070 157.255 ;
    END
  END addr_r1[1]
  PIN addr_r1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.005 0.070 159.075 ;
    END
  END addr_r1[2]
  PIN addr_r1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.825 0.070 160.895 ;
    END
  END addr_r1[3]
  PIN addr_r1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.645 0.070 162.715 ;
    END
  END addr_r1[4]
  PIN addr_r1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.465 0.070 164.535 ;
    END
  END addr_r1[5]
  PIN addr_r2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.865 0.070 165.935 ;
    END
  END addr_r2[0]
  PIN addr_r2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.685 0.070 167.755 ;
    END
  END addr_r2[1]
  PIN addr_r2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.505 0.070 169.575 ;
    END
  END addr_r2[2]
  PIN addr_r2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.325 0.070 171.395 ;
    END
  END addr_r2[3]
  PIN addr_r2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.145 0.070 173.215 ;
    END
  END addr_r2[4]
  PIN addr_r2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.965 0.070 175.035 ;
    END
  END addr_r2[5]
  PIN we_in_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.365 0.070 176.435 ;
    END
  END we_in_w1
  PIN ce_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.345 0.070 177.415 ;
    END
  END ce_w1
  PIN ce_r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.745 0.070 178.815 ;
    END
  END ce_r1
  PIN ce_r2
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.565 0.070 180.635 ;
    END
  END ce_r2
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.965 0.070 182.035 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 133.000 ;
      RECT 3.500 1.400 3.780 133.000 ;
      RECT 5.740 1.400 6.020 133.000 ;
      RECT 7.980 1.400 8.260 133.000 ;
      RECT 10.220 1.400 10.500 133.000 ;
      RECT 12.460 1.400 12.740 133.000 ;
      RECT 14.700 1.400 14.980 133.000 ;
      RECT 16.940 1.400 17.220 133.000 ;
      RECT 19.180 1.400 19.460 133.000 ;
      RECT 21.420 1.400 21.700 133.000 ;
      RECT 23.660 1.400 23.940 133.000 ;
      RECT 25.900 1.400 26.180 133.000 ;
      RECT 28.140 1.400 28.420 133.000 ;
      RECT 30.380 1.400 30.660 133.000 ;
      RECT 32.620 1.400 32.900 133.000 ;
      RECT 34.860 1.400 35.140 133.000 ;
      RECT 37.100 1.400 37.380 133.000 ;
      RECT 39.340 1.400 39.620 133.000 ;
      RECT 41.580 1.400 41.860 133.000 ;
      RECT 43.820 1.400 44.100 133.000 ;
      RECT 46.060 1.400 46.340 133.000 ;
      RECT 48.300 1.400 48.580 133.000 ;
      RECT 50.540 1.400 50.820 133.000 ;
      RECT 52.780 1.400 53.060 133.000 ;
      RECT 55.020 1.400 55.300 133.000 ;
      RECT 57.260 1.400 57.540 133.000 ;
      RECT 59.500 1.400 59.780 133.000 ;
      RECT 61.740 1.400 62.020 133.000 ;
      RECT 63.980 1.400 64.260 133.000 ;
      RECT 66.220 1.400 66.500 133.000 ;
      RECT 68.460 1.400 68.740 133.000 ;
      RECT 70.700 1.400 70.980 133.000 ;
      RECT 72.940 1.400 73.220 133.000 ;
      RECT 75.180 1.400 75.460 133.000 ;
      RECT 77.420 1.400 77.700 133.000 ;
      RECT 79.660 1.400 79.940 133.000 ;
      RECT 81.900 1.400 82.180 133.000 ;
      RECT 84.140 1.400 84.420 133.000 ;
      RECT 86.380 1.400 86.660 133.000 ;
      RECT 88.620 1.400 88.900 133.000 ;
      RECT 90.860 1.400 91.140 133.000 ;
      RECT 93.100 1.400 93.380 133.000 ;
      RECT 95.340 1.400 95.620 133.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 133.000 ;
      RECT 4.620 1.400 4.900 133.000 ;
      RECT 6.860 1.400 7.140 133.000 ;
      RECT 9.100 1.400 9.380 133.000 ;
      RECT 11.340 1.400 11.620 133.000 ;
      RECT 13.580 1.400 13.860 133.000 ;
      RECT 15.820 1.400 16.100 133.000 ;
      RECT 18.060 1.400 18.340 133.000 ;
      RECT 20.300 1.400 20.580 133.000 ;
      RECT 22.540 1.400 22.820 133.000 ;
      RECT 24.780 1.400 25.060 133.000 ;
      RECT 27.020 1.400 27.300 133.000 ;
      RECT 29.260 1.400 29.540 133.000 ;
      RECT 31.500 1.400 31.780 133.000 ;
      RECT 33.740 1.400 34.020 133.000 ;
      RECT 35.980 1.400 36.260 133.000 ;
      RECT 38.220 1.400 38.500 133.000 ;
      RECT 40.460 1.400 40.740 133.000 ;
      RECT 42.700 1.400 42.980 133.000 ;
      RECT 44.940 1.400 45.220 133.000 ;
      RECT 47.180 1.400 47.460 133.000 ;
      RECT 49.420 1.400 49.700 133.000 ;
      RECT 51.660 1.400 51.940 133.000 ;
      RECT 53.900 1.400 54.180 133.000 ;
      RECT 56.140 1.400 56.420 133.000 ;
      RECT 58.380 1.400 58.660 133.000 ;
      RECT 60.620 1.400 60.900 133.000 ;
      RECT 62.860 1.400 63.140 133.000 ;
      RECT 65.100 1.400 65.380 133.000 ;
      RECT 67.340 1.400 67.620 133.000 ;
      RECT 69.580 1.400 69.860 133.000 ;
      RECT 71.820 1.400 72.100 133.000 ;
      RECT 74.060 1.400 74.340 133.000 ;
      RECT 76.300 1.400 76.580 133.000 ;
      RECT 78.540 1.400 78.820 133.000 ;
      RECT 80.780 1.400 81.060 133.000 ;
      RECT 83.020 1.400 83.300 133.000 ;
      RECT 85.260 1.400 85.540 133.000 ;
      RECT 87.500 1.400 87.780 133.000 ;
      RECT 89.740 1.400 90.020 133.000 ;
      RECT 91.980 1.400 92.260 133.000 ;
      RECT 94.220 1.400 94.500 133.000 ;
      RECT 96.460 1.400 96.740 133.000 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 98.990 134.400 ;
    LAYER metal2 ;
    RECT 0 0 98.990 134.400 ;
    LAYER metal3 ;
    RECT 0.070 0 98.990 134.400 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 3.185 ;
    RECT 0 3.255 0.070 5.005 ;
    RECT 0 5.075 0.070 6.825 ;
    RECT 0 6.895 0.070 8.645 ;
    RECT 0 8.715 0.070 10.465 ;
    RECT 0 10.535 0.070 12.285 ;
    RECT 0 12.355 0.070 14.105 ;
    RECT 0 14.175 0.070 15.925 ;
    RECT 0 15.995 0.070 17.745 ;
    RECT 0 17.815 0.070 19.565 ;
    RECT 0 19.635 0.070 21.385 ;
    RECT 0 21.455 0.070 23.205 ;
    RECT 0 23.275 0.070 25.025 ;
    RECT 0 25.095 0.070 26.845 ;
    RECT 0 26.915 0.070 28.665 ;
    RECT 0 28.735 0.070 30.485 ;
    RECT 0 30.555 0.070 32.305 ;
    RECT 0 32.375 0.070 34.125 ;
    RECT 0 34.195 0.070 35.945 ;
    RECT 0 36.015 0.070 37.345 ;
    RECT 0 37.415 0.070 39.165 ;
    RECT 0 39.235 0.070 40.985 ;
    RECT 0 41.055 0.070 42.805 ;
    RECT 0 42.875 0.070 44.625 ;
    RECT 0 44.695 0.070 46.445 ;
    RECT 0 46.515 0.070 48.265 ;
    RECT 0 48.335 0.070 50.085 ;
    RECT 0 50.155 0.070 51.905 ;
    RECT 0 51.975 0.070 53.725 ;
    RECT 0 53.795 0.070 55.545 ;
    RECT 0 55.615 0.070 57.365 ;
    RECT 0 57.435 0.070 59.185 ;
    RECT 0 59.255 0.070 61.005 ;
    RECT 0 61.075 0.070 62.825 ;
    RECT 0 62.895 0.070 64.645 ;
    RECT 0 64.715 0.070 66.465 ;
    RECT 0 66.535 0.070 68.285 ;
    RECT 0 68.355 0.070 70.105 ;
    RECT 0 70.175 0.070 71.925 ;
    RECT 0 71.995 0.070 73.325 ;
    RECT 0 73.395 0.070 75.145 ;
    RECT 0 75.215 0.070 76.965 ;
    RECT 0 77.035 0.070 78.785 ;
    RECT 0 78.855 0.070 80.605 ;
    RECT 0 80.675 0.070 82.425 ;
    RECT 0 82.495 0.070 84.245 ;
    RECT 0 84.315 0.070 86.065 ;
    RECT 0 86.135 0.070 87.885 ;
    RECT 0 87.955 0.070 89.705 ;
    RECT 0 89.775 0.070 91.525 ;
    RECT 0 91.595 0.070 93.345 ;
    RECT 0 93.415 0.070 95.165 ;
    RECT 0 95.235 0.070 96.985 ;
    RECT 0 97.055 0.070 98.805 ;
    RECT 0 98.875 0.070 100.625 ;
    RECT 0 100.695 0.070 102.445 ;
    RECT 0 102.515 0.070 104.265 ;
    RECT 0 104.335 0.070 106.085 ;
    RECT 0 106.155 0.070 107.905 ;
    RECT 0 107.975 0.070 109.305 ;
    RECT 0 109.375 0.070 111.125 ;
    RECT 0 111.195 0.070 112.945 ;
    RECT 0 113.015 0.070 114.765 ;
    RECT 0 114.835 0.070 116.585 ;
    RECT 0 116.655 0.070 118.405 ;
    RECT 0 118.475 0.070 119.805 ;
    RECT 0 119.875 0.070 121.625 ;
    RECT 0 121.695 0.070 123.445 ;
    RECT 0 123.515 0.070 134.400 ;
    LAYER metal4 ;
    RECT 0 0 98.990 1.400 ;
    RECT 0 133.000 98.990 134.400 ;
    RECT 0.000 1.400 1.260 133.000 ;
    RECT 1.540 1.400 2.380 133.000 ;
    RECT 2.660 1.400 3.500 133.000 ;
    RECT 3.780 1.400 4.620 133.000 ;
    RECT 4.900 1.400 5.740 133.000 ;
    RECT 6.020 1.400 6.860 133.000 ;
    RECT 7.140 1.400 7.980 133.000 ;
    RECT 8.260 1.400 9.100 133.000 ;
    RECT 9.380 1.400 10.220 133.000 ;
    RECT 10.500 1.400 11.340 133.000 ;
    RECT 11.620 1.400 12.460 133.000 ;
    RECT 12.740 1.400 13.580 133.000 ;
    RECT 13.860 1.400 14.700 133.000 ;
    RECT 14.980 1.400 15.820 133.000 ;
    RECT 16.100 1.400 16.940 133.000 ;
    RECT 17.220 1.400 18.060 133.000 ;
    RECT 18.340 1.400 19.180 133.000 ;
    RECT 19.460 1.400 20.300 133.000 ;
    RECT 20.580 1.400 21.420 133.000 ;
    RECT 21.700 1.400 22.540 133.000 ;
    RECT 22.820 1.400 23.660 133.000 ;
    RECT 23.940 1.400 24.780 133.000 ;
    RECT 25.060 1.400 25.900 133.000 ;
    RECT 26.180 1.400 27.020 133.000 ;
    RECT 27.300 1.400 28.140 133.000 ;
    RECT 28.420 1.400 29.260 133.000 ;
    RECT 29.540 1.400 30.380 133.000 ;
    RECT 30.660 1.400 31.500 133.000 ;
    RECT 31.780 1.400 32.620 133.000 ;
    RECT 32.900 1.400 33.740 133.000 ;
    RECT 34.020 1.400 34.860 133.000 ;
    RECT 35.140 1.400 35.980 133.000 ;
    RECT 36.260 1.400 37.100 133.000 ;
    RECT 37.380 1.400 38.220 133.000 ;
    RECT 38.500 1.400 39.340 133.000 ;
    RECT 39.620 1.400 40.460 133.000 ;
    RECT 40.740 1.400 41.580 133.000 ;
    RECT 41.860 1.400 42.700 133.000 ;
    RECT 42.980 1.400 43.820 133.000 ;
    RECT 44.100 1.400 44.940 133.000 ;
    RECT 45.220 1.400 46.060 133.000 ;
    RECT 46.340 1.400 47.180 133.000 ;
    RECT 47.460 1.400 48.300 133.000 ;
    RECT 48.580 1.400 49.420 133.000 ;
    RECT 49.700 1.400 50.540 133.000 ;
    RECT 50.820 1.400 51.660 133.000 ;
    RECT 51.940 1.400 52.780 133.000 ;
    RECT 53.060 1.400 53.900 133.000 ;
    RECT 54.180 1.400 55.020 133.000 ;
    RECT 55.300 1.400 56.140 133.000 ;
    RECT 56.420 1.400 57.260 133.000 ;
    RECT 57.540 1.400 58.380 133.000 ;
    RECT 58.660 1.400 59.500 133.000 ;
    RECT 59.780 1.400 60.620 133.000 ;
    RECT 60.900 1.400 61.740 133.000 ;
    RECT 62.020 1.400 62.860 133.000 ;
    RECT 63.140 1.400 63.980 133.000 ;
    RECT 64.260 1.400 65.100 133.000 ;
    RECT 65.380 1.400 66.220 133.000 ;
    RECT 66.500 1.400 67.340 133.000 ;
    RECT 67.620 1.400 68.460 133.000 ;
    RECT 68.740 1.400 69.580 133.000 ;
    RECT 69.860 1.400 70.700 133.000 ;
    RECT 70.980 1.400 71.820 133.000 ;
    RECT 72.100 1.400 72.940 133.000 ;
    RECT 73.220 1.400 74.060 133.000 ;
    RECT 74.340 1.400 75.180 133.000 ;
    RECT 75.460 1.400 76.300 133.000 ;
    RECT 76.580 1.400 77.420 133.000 ;
    RECT 77.700 1.400 78.540 133.000 ;
    RECT 78.820 1.400 79.660 133.000 ;
    RECT 79.940 1.400 80.780 133.000 ;
    RECT 81.060 1.400 81.900 133.000 ;
    RECT 82.180 1.400 83.020 133.000 ;
    RECT 83.300 1.400 84.140 133.000 ;
    RECT 84.420 1.400 85.260 133.000 ;
    RECT 85.540 1.400 86.380 133.000 ;
    RECT 86.660 1.400 87.500 133.000 ;
    RECT 87.780 1.400 88.620 133.000 ;
    RECT 88.900 1.400 89.740 133.000 ;
    RECT 90.020 1.400 90.860 133.000 ;
    RECT 91.140 1.400 91.980 133.000 ;
    RECT 92.260 1.400 93.100 133.000 ;
    RECT 93.380 1.400 94.220 133.000 ;
    RECT 94.500 1.400 95.340 133.000 ;
    RECT 95.620 1.400 96.460 133.000 ;
    RECT 96.740 1.400 98.990 133.000 ;
    LAYER OVERLAP ;
    RECT 0 0 98.990 134.400 ;
  END
END fakeram_20x64_2r1w

END LIBRARY
