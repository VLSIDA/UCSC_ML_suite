VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_32x1024_2r1w
  FOREIGN sram_32x1024_2r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 209.000 BY 642.600 ;
  CLASS BLOCK ;
  PIN w_mask_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 -0.875 0.070 -0.805 ;
    END
  END w_mask_w1[0]
  PIN w_mask_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.865 0.070 4.935 ;
    END
  END w_mask_w1[1]
  PIN w_mask_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_w1[2]
  PIN w_mask_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_w1[3]
  PIN w_mask_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.085 0.070 22.155 ;
    END
  END w_mask_w1[4]
  PIN w_mask_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.825 0.070 27.895 ;
    END
  END w_mask_w1[5]
  PIN w_mask_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END w_mask_w1[6]
  PIN w_mask_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.305 0.070 39.375 ;
    END
  END w_mask_w1[7]
  PIN w_mask_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END w_mask_w1[8]
  PIN w_mask_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END w_mask_w1[9]
  PIN w_mask_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.525 0.070 56.595 ;
    END
  END w_mask_w1[10]
  PIN w_mask_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.265 0.070 62.335 ;
    END
  END w_mask_w1[11]
  PIN w_mask_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END w_mask_w1[12]
  PIN w_mask_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.745 0.070 73.815 ;
    END
  END w_mask_w1[13]
  PIN w_mask_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.485 0.070 79.555 ;
    END
  END w_mask_w1[14]
  PIN w_mask_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END w_mask_w1[15]
  PIN w_mask_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.965 0.070 91.035 ;
    END
  END w_mask_w1[16]
  PIN w_mask_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.705 0.070 96.775 ;
    END
  END w_mask_w1[17]
  PIN w_mask_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.445 0.070 102.515 ;
    END
  END w_mask_w1[18]
  PIN w_mask_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.185 0.070 108.255 ;
    END
  END w_mask_w1[19]
  PIN w_mask_w1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.925 0.070 113.995 ;
    END
  END w_mask_w1[20]
  PIN w_mask_w1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.665 0.070 119.735 ;
    END
  END w_mask_w1[21]
  PIN w_mask_w1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.405 0.070 125.475 ;
    END
  END w_mask_w1[22]
  PIN w_mask_w1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.145 0.070 131.215 ;
    END
  END w_mask_w1[23]
  PIN w_mask_w1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.885 0.070 136.955 ;
    END
  END w_mask_w1[24]
  PIN w_mask_w1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.625 0.070 142.695 ;
    END
  END w_mask_w1[25]
  PIN w_mask_w1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.365 0.070 148.435 ;
    END
  END w_mask_w1[26]
  PIN w_mask_w1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.105 0.070 154.175 ;
    END
  END w_mask_w1[27]
  PIN w_mask_w1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.845 0.070 159.915 ;
    END
  END w_mask_w1[28]
  PIN w_mask_w1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.585 0.070 165.655 ;
    END
  END w_mask_w1[29]
  PIN w_mask_w1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.325 0.070 171.395 ;
    END
  END w_mask_w1[30]
  PIN w_mask_w1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.065 0.070 177.135 ;
    END
  END w_mask_w1[31]
  PIN rd_out_r1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.565 0.070 180.635 ;
    END
  END rd_out_r1[0]
  PIN rd_out_r1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.305 0.070 186.375 ;
    END
  END rd_out_r1[1]
  PIN rd_out_r1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.045 0.070 192.115 ;
    END
  END rd_out_r1[2]
  PIN rd_out_r1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.785 0.070 197.855 ;
    END
  END rd_out_r1[3]
  PIN rd_out_r1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.525 0.070 203.595 ;
    END
  END rd_out_r1[4]
  PIN rd_out_r1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.265 0.070 209.335 ;
    END
  END rd_out_r1[5]
  PIN rd_out_r1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.005 0.070 215.075 ;
    END
  END rd_out_r1[6]
  PIN rd_out_r1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.745 0.070 220.815 ;
    END
  END rd_out_r1[7]
  PIN rd_out_r1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.485 0.070 226.555 ;
    END
  END rd_out_r1[8]
  PIN rd_out_r1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.225 0.070 232.295 ;
    END
  END rd_out_r1[9]
  PIN rd_out_r1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.965 0.070 238.035 ;
    END
  END rd_out_r1[10]
  PIN rd_out_r1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.705 0.070 243.775 ;
    END
  END rd_out_r1[11]
  PIN rd_out_r1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.445 0.070 249.515 ;
    END
  END rd_out_r1[12]
  PIN rd_out_r1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.185 0.070 255.255 ;
    END
  END rd_out_r1[13]
  PIN rd_out_r1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.925 0.070 260.995 ;
    END
  END rd_out_r1[14]
  PIN rd_out_r1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.665 0.070 266.735 ;
    END
  END rd_out_r1[15]
  PIN rd_out_r1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.405 0.070 272.475 ;
    END
  END rd_out_r1[16]
  PIN rd_out_r1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.145 0.070 278.215 ;
    END
  END rd_out_r1[17]
  PIN rd_out_r1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.885 0.070 283.955 ;
    END
  END rd_out_r1[18]
  PIN rd_out_r1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.625 0.070 289.695 ;
    END
  END rd_out_r1[19]
  PIN rd_out_r1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.365 0.070 295.435 ;
    END
  END rd_out_r1[20]
  PIN rd_out_r1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.105 0.070 301.175 ;
    END
  END rd_out_r1[21]
  PIN rd_out_r1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.845 0.070 306.915 ;
    END
  END rd_out_r1[22]
  PIN rd_out_r1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.585 0.070 312.655 ;
    END
  END rd_out_r1[23]
  PIN rd_out_r1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.325 0.070 318.395 ;
    END
  END rd_out_r1[24]
  PIN rd_out_r1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.065 0.070 324.135 ;
    END
  END rd_out_r1[25]
  PIN rd_out_r1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.805 0.070 329.875 ;
    END
  END rd_out_r1[26]
  PIN rd_out_r1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.545 0.070 335.615 ;
    END
  END rd_out_r1[27]
  PIN rd_out_r1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.285 0.070 341.355 ;
    END
  END rd_out_r1[28]
  PIN rd_out_r1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.025 0.070 347.095 ;
    END
  END rd_out_r1[29]
  PIN rd_out_r1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.765 0.070 352.835 ;
    END
  END rd_out_r1[30]
  PIN rd_out_r1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.505 0.070 358.575 ;
    END
  END rd_out_r1[31]
  PIN rd_out_r2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.005 0.070 362.075 ;
    END
  END rd_out_r2[0]
  PIN rd_out_r2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.745 0.070 367.815 ;
    END
  END rd_out_r2[1]
  PIN rd_out_r2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.485 0.070 373.555 ;
    END
  END rd_out_r2[2]
  PIN rd_out_r2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.225 0.070 379.295 ;
    END
  END rd_out_r2[3]
  PIN rd_out_r2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.965 0.070 385.035 ;
    END
  END rd_out_r2[4]
  PIN rd_out_r2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.705 0.070 390.775 ;
    END
  END rd_out_r2[5]
  PIN rd_out_r2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.445 0.070 396.515 ;
    END
  END rd_out_r2[6]
  PIN rd_out_r2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 402.185 0.070 402.255 ;
    END
  END rd_out_r2[7]
  PIN rd_out_r2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 407.925 0.070 407.995 ;
    END
  END rd_out_r2[8]
  PIN rd_out_r2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 413.665 0.070 413.735 ;
    END
  END rd_out_r2[9]
  PIN rd_out_r2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 419.405 0.070 419.475 ;
    END
  END rd_out_r2[10]
  PIN rd_out_r2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 425.145 0.070 425.215 ;
    END
  END rd_out_r2[11]
  PIN rd_out_r2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 430.885 0.070 430.955 ;
    END
  END rd_out_r2[12]
  PIN rd_out_r2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 436.625 0.070 436.695 ;
    END
  END rd_out_r2[13]
  PIN rd_out_r2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 442.365 0.070 442.435 ;
    END
  END rd_out_r2[14]
  PIN rd_out_r2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 448.105 0.070 448.175 ;
    END
  END rd_out_r2[15]
  PIN rd_out_r2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 453.845 0.070 453.915 ;
    END
  END rd_out_r2[16]
  PIN rd_out_r2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 459.585 0.070 459.655 ;
    END
  END rd_out_r2[17]
  PIN rd_out_r2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 465.325 0.070 465.395 ;
    END
  END rd_out_r2[18]
  PIN rd_out_r2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 471.065 0.070 471.135 ;
    END
  END rd_out_r2[19]
  PIN rd_out_r2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 476.805 0.070 476.875 ;
    END
  END rd_out_r2[20]
  PIN rd_out_r2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 482.545 0.070 482.615 ;
    END
  END rd_out_r2[21]
  PIN rd_out_r2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 488.285 0.070 488.355 ;
    END
  END rd_out_r2[22]
  PIN rd_out_r2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 494.025 0.070 494.095 ;
    END
  END rd_out_r2[23]
  PIN rd_out_r2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 499.765 0.070 499.835 ;
    END
  END rd_out_r2[24]
  PIN rd_out_r2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.505 0.070 505.575 ;
    END
  END rd_out_r2[25]
  PIN rd_out_r2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 511.245 0.070 511.315 ;
    END
  END rd_out_r2[26]
  PIN rd_out_r2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.985 0.070 517.055 ;
    END
  END rd_out_r2[27]
  PIN rd_out_r2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.725 0.070 522.795 ;
    END
  END rd_out_r2[28]
  PIN rd_out_r2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.465 0.070 528.535 ;
    END
  END rd_out_r2[29]
  PIN rd_out_r2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.205 0.070 534.275 ;
    END
  END rd_out_r2[30]
  PIN rd_out_r2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.945 0.070 540.015 ;
    END
  END rd_out_r2[31]
  PIN wd_in_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.445 0.070 543.515 ;
    END
  END wd_in_w1[0]
  PIN wd_in_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.185 0.070 549.255 ;
    END
  END wd_in_w1[1]
  PIN wd_in_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.925 0.070 554.995 ;
    END
  END wd_in_w1[2]
  PIN wd_in_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.665 0.070 560.735 ;
    END
  END wd_in_w1[3]
  PIN wd_in_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.405 0.070 566.475 ;
    END
  END wd_in_w1[4]
  PIN wd_in_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.145 0.070 572.215 ;
    END
  END wd_in_w1[5]
  PIN wd_in_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.885 0.070 577.955 ;
    END
  END wd_in_w1[6]
  PIN wd_in_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.625 0.070 583.695 ;
    END
  END wd_in_w1[7]
  PIN wd_in_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.365 0.070 589.435 ;
    END
  END wd_in_w1[8]
  PIN wd_in_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.105 0.070 595.175 ;
    END
  END wd_in_w1[9]
  PIN wd_in_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.845 0.070 600.915 ;
    END
  END wd_in_w1[10]
  PIN wd_in_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.585 0.070 606.655 ;
    END
  END wd_in_w1[11]
  PIN wd_in_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.325 0.070 612.395 ;
    END
  END wd_in_w1[12]
  PIN wd_in_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.065 0.070 618.135 ;
    END
  END wd_in_w1[13]
  PIN wd_in_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.805 0.070 623.875 ;
    END
  END wd_in_w1[14]
  PIN wd_in_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 629.545 0.070 629.615 ;
    END
  END wd_in_w1[15]
  PIN wd_in_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.285 0.070 635.355 ;
    END
  END wd_in_w1[16]
  PIN wd_in_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.025 0.070 641.095 ;
    END
  END wd_in_w1[17]
  PIN wd_in_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.765 0.070 646.835 ;
    END
  END wd_in_w1[18]
  PIN wd_in_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.505 0.070 652.575 ;
    END
  END wd_in_w1[19]
  PIN wd_in_w1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.245 0.070 658.315 ;
    END
  END wd_in_w1[20]
  PIN wd_in_w1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.985 0.070 664.055 ;
    END
  END wd_in_w1[21]
  PIN wd_in_w1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.725 0.070 669.795 ;
    END
  END wd_in_w1[22]
  PIN wd_in_w1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.465 0.070 675.535 ;
    END
  END wd_in_w1[23]
  PIN wd_in_w1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.205 0.070 681.275 ;
    END
  END wd_in_w1[24]
  PIN wd_in_w1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 686.945 0.070 687.015 ;
    END
  END wd_in_w1[25]
  PIN wd_in_w1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.685 0.070 692.755 ;
    END
  END wd_in_w1[26]
  PIN wd_in_w1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.425 0.070 698.495 ;
    END
  END wd_in_w1[27]
  PIN wd_in_w1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.165 0.070 704.235 ;
    END
  END wd_in_w1[28]
  PIN wd_in_w1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.905 0.070 709.975 ;
    END
  END wd_in_w1[29]
  PIN wd_in_w1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.645 0.070 715.715 ;
    END
  END wd_in_w1[30]
  PIN wd_in_w1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.385 0.070 721.455 ;
    END
  END wd_in_w1[31]
  PIN addr_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.885 0.070 724.955 ;
    END
  END addr_w1[0]
  PIN addr_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.625 0.070 730.695 ;
    END
  END addr_w1[1]
  PIN addr_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 736.365 0.070 736.435 ;
    END
  END addr_w1[2]
  PIN addr_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 742.105 0.070 742.175 ;
    END
  END addr_w1[3]
  PIN addr_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.845 0.070 747.915 ;
    END
  END addr_w1[4]
  PIN addr_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 753.585 0.070 753.655 ;
    END
  END addr_w1[5]
  PIN addr_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.325 0.070 759.395 ;
    END
  END addr_w1[6]
  PIN addr_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 765.065 0.070 765.135 ;
    END
  END addr_w1[7]
  PIN addr_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 770.805 0.070 770.875 ;
    END
  END addr_w1[8]
  PIN addr_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 776.545 0.070 776.615 ;
    END
  END addr_w1[9]
  PIN addr_r1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 780.045 0.070 780.115 ;
    END
  END addr_r1[0]
  PIN addr_r1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 785.785 0.070 785.855 ;
    END
  END addr_r1[1]
  PIN addr_r1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 791.525 0.070 791.595 ;
    END
  END addr_r1[2]
  PIN addr_r1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 797.265 0.070 797.335 ;
    END
  END addr_r1[3]
  PIN addr_r1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 803.005 0.070 803.075 ;
    END
  END addr_r1[4]
  PIN addr_r1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 808.745 0.070 808.815 ;
    END
  END addr_r1[5]
  PIN addr_r1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 814.485 0.070 814.555 ;
    END
  END addr_r1[6]
  PIN addr_r1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 820.225 0.070 820.295 ;
    END
  END addr_r1[7]
  PIN addr_r1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 825.965 0.070 826.035 ;
    END
  END addr_r1[8]
  PIN addr_r1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.705 0.070 831.775 ;
    END
  END addr_r1[9]
  PIN addr_r2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 835.205 0.070 835.275 ;
    END
  END addr_r2[0]
  PIN addr_r2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 840.945 0.070 841.015 ;
    END
  END addr_r2[1]
  PIN addr_r2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 846.685 0.070 846.755 ;
    END
  END addr_r2[2]
  PIN addr_r2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.425 0.070 852.495 ;
    END
  END addr_r2[3]
  PIN addr_r2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 858.165 0.070 858.235 ;
    END
  END addr_r2[4]
  PIN addr_r2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 863.905 0.070 863.975 ;
    END
  END addr_r2[5]
  PIN addr_r2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 869.645 0.070 869.715 ;
    END
  END addr_r2[6]
  PIN addr_r2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 875.385 0.070 875.455 ;
    END
  END addr_r2[7]
  PIN addr_r2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 881.125 0.070 881.195 ;
    END
  END addr_r2[8]
  PIN addr_r2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 886.865 0.070 886.935 ;
    END
  END addr_r2[9]
  PIN we_in_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 890.365 0.070 890.435 ;
    END
  END we_in_w1
  PIN ce_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 891.625 0.070 891.695 ;
    END
  END ce_w1
  PIN ce_r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 895.125 0.070 895.195 ;
    END
  END ce_r1
  PIN ce_r2
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 900.865 0.070 900.935 ;
    END
  END ce_r2
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 904.365 0.070 904.435 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 641.200 ;
      RECT 3.500 1.400 3.780 641.200 ;
      RECT 5.740 1.400 6.020 641.200 ;
      RECT 7.980 1.400 8.260 641.200 ;
      RECT 10.220 1.400 10.500 641.200 ;
      RECT 12.460 1.400 12.740 641.200 ;
      RECT 14.700 1.400 14.980 641.200 ;
      RECT 16.940 1.400 17.220 641.200 ;
      RECT 19.180 1.400 19.460 641.200 ;
      RECT 21.420 1.400 21.700 641.200 ;
      RECT 23.660 1.400 23.940 641.200 ;
      RECT 25.900 1.400 26.180 641.200 ;
      RECT 28.140 1.400 28.420 641.200 ;
      RECT 30.380 1.400 30.660 641.200 ;
      RECT 32.620 1.400 32.900 641.200 ;
      RECT 34.860 1.400 35.140 641.200 ;
      RECT 37.100 1.400 37.380 641.200 ;
      RECT 39.340 1.400 39.620 641.200 ;
      RECT 41.580 1.400 41.860 641.200 ;
      RECT 43.820 1.400 44.100 641.200 ;
      RECT 46.060 1.400 46.340 641.200 ;
      RECT 48.300 1.400 48.580 641.200 ;
      RECT 50.540 1.400 50.820 641.200 ;
      RECT 52.780 1.400 53.060 641.200 ;
      RECT 55.020 1.400 55.300 641.200 ;
      RECT 57.260 1.400 57.540 641.200 ;
      RECT 59.500 1.400 59.780 641.200 ;
      RECT 61.740 1.400 62.020 641.200 ;
      RECT 63.980 1.400 64.260 641.200 ;
      RECT 66.220 1.400 66.500 641.200 ;
      RECT 68.460 1.400 68.740 641.200 ;
      RECT 70.700 1.400 70.980 641.200 ;
      RECT 72.940 1.400 73.220 641.200 ;
      RECT 75.180 1.400 75.460 641.200 ;
      RECT 77.420 1.400 77.700 641.200 ;
      RECT 79.660 1.400 79.940 641.200 ;
      RECT 81.900 1.400 82.180 641.200 ;
      RECT 84.140 1.400 84.420 641.200 ;
      RECT 86.380 1.400 86.660 641.200 ;
      RECT 88.620 1.400 88.900 641.200 ;
      RECT 90.860 1.400 91.140 641.200 ;
      RECT 93.100 1.400 93.380 641.200 ;
      RECT 95.340 1.400 95.620 641.200 ;
      RECT 97.580 1.400 97.860 641.200 ;
      RECT 99.820 1.400 100.100 641.200 ;
      RECT 102.060 1.400 102.340 641.200 ;
      RECT 104.300 1.400 104.580 641.200 ;
      RECT 106.540 1.400 106.820 641.200 ;
      RECT 108.780 1.400 109.060 641.200 ;
      RECT 111.020 1.400 111.300 641.200 ;
      RECT 113.260 1.400 113.540 641.200 ;
      RECT 115.500 1.400 115.780 641.200 ;
      RECT 117.740 1.400 118.020 641.200 ;
      RECT 119.980 1.400 120.260 641.200 ;
      RECT 122.220 1.400 122.500 641.200 ;
      RECT 124.460 1.400 124.740 641.200 ;
      RECT 126.700 1.400 126.980 641.200 ;
      RECT 128.940 1.400 129.220 641.200 ;
      RECT 131.180 1.400 131.460 641.200 ;
      RECT 133.420 1.400 133.700 641.200 ;
      RECT 135.660 1.400 135.940 641.200 ;
      RECT 137.900 1.400 138.180 641.200 ;
      RECT 140.140 1.400 140.420 641.200 ;
      RECT 142.380 1.400 142.660 641.200 ;
      RECT 144.620 1.400 144.900 641.200 ;
      RECT 146.860 1.400 147.140 641.200 ;
      RECT 149.100 1.400 149.380 641.200 ;
      RECT 151.340 1.400 151.620 641.200 ;
      RECT 153.580 1.400 153.860 641.200 ;
      RECT 155.820 1.400 156.100 641.200 ;
      RECT 158.060 1.400 158.340 641.200 ;
      RECT 160.300 1.400 160.580 641.200 ;
      RECT 162.540 1.400 162.820 641.200 ;
      RECT 164.780 1.400 165.060 641.200 ;
      RECT 167.020 1.400 167.300 641.200 ;
      RECT 169.260 1.400 169.540 641.200 ;
      RECT 171.500 1.400 171.780 641.200 ;
      RECT 173.740 1.400 174.020 641.200 ;
      RECT 175.980 1.400 176.260 641.200 ;
      RECT 178.220 1.400 178.500 641.200 ;
      RECT 180.460 1.400 180.740 641.200 ;
      RECT 182.700 1.400 182.980 641.200 ;
      RECT 184.940 1.400 185.220 641.200 ;
      RECT 187.180 1.400 187.460 641.200 ;
      RECT 189.420 1.400 189.700 641.200 ;
      RECT 191.660 1.400 191.940 641.200 ;
      RECT 193.900 1.400 194.180 641.200 ;
      RECT 196.140 1.400 196.420 641.200 ;
      RECT 198.380 1.400 198.660 641.200 ;
      RECT 200.620 1.400 200.900 641.200 ;
      RECT 202.860 1.400 203.140 641.200 ;
      RECT 205.100 1.400 205.380 641.200 ;
      RECT 207.340 1.400 207.620 641.200 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 641.200 ;
      RECT 4.620 1.400 4.900 641.200 ;
      RECT 6.860 1.400 7.140 641.200 ;
      RECT 9.100 1.400 9.380 641.200 ;
      RECT 11.340 1.400 11.620 641.200 ;
      RECT 13.580 1.400 13.860 641.200 ;
      RECT 15.820 1.400 16.100 641.200 ;
      RECT 18.060 1.400 18.340 641.200 ;
      RECT 20.300 1.400 20.580 641.200 ;
      RECT 22.540 1.400 22.820 641.200 ;
      RECT 24.780 1.400 25.060 641.200 ;
      RECT 27.020 1.400 27.300 641.200 ;
      RECT 29.260 1.400 29.540 641.200 ;
      RECT 31.500 1.400 31.780 641.200 ;
      RECT 33.740 1.400 34.020 641.200 ;
      RECT 35.980 1.400 36.260 641.200 ;
      RECT 38.220 1.400 38.500 641.200 ;
      RECT 40.460 1.400 40.740 641.200 ;
      RECT 42.700 1.400 42.980 641.200 ;
      RECT 44.940 1.400 45.220 641.200 ;
      RECT 47.180 1.400 47.460 641.200 ;
      RECT 49.420 1.400 49.700 641.200 ;
      RECT 51.660 1.400 51.940 641.200 ;
      RECT 53.900 1.400 54.180 641.200 ;
      RECT 56.140 1.400 56.420 641.200 ;
      RECT 58.380 1.400 58.660 641.200 ;
      RECT 60.620 1.400 60.900 641.200 ;
      RECT 62.860 1.400 63.140 641.200 ;
      RECT 65.100 1.400 65.380 641.200 ;
      RECT 67.340 1.400 67.620 641.200 ;
      RECT 69.580 1.400 69.860 641.200 ;
      RECT 71.820 1.400 72.100 641.200 ;
      RECT 74.060 1.400 74.340 641.200 ;
      RECT 76.300 1.400 76.580 641.200 ;
      RECT 78.540 1.400 78.820 641.200 ;
      RECT 80.780 1.400 81.060 641.200 ;
      RECT 83.020 1.400 83.300 641.200 ;
      RECT 85.260 1.400 85.540 641.200 ;
      RECT 87.500 1.400 87.780 641.200 ;
      RECT 89.740 1.400 90.020 641.200 ;
      RECT 91.980 1.400 92.260 641.200 ;
      RECT 94.220 1.400 94.500 641.200 ;
      RECT 96.460 1.400 96.740 641.200 ;
      RECT 98.700 1.400 98.980 641.200 ;
      RECT 100.940 1.400 101.220 641.200 ;
      RECT 103.180 1.400 103.460 641.200 ;
      RECT 105.420 1.400 105.700 641.200 ;
      RECT 107.660 1.400 107.940 641.200 ;
      RECT 109.900 1.400 110.180 641.200 ;
      RECT 112.140 1.400 112.420 641.200 ;
      RECT 114.380 1.400 114.660 641.200 ;
      RECT 116.620 1.400 116.900 641.200 ;
      RECT 118.860 1.400 119.140 641.200 ;
      RECT 121.100 1.400 121.380 641.200 ;
      RECT 123.340 1.400 123.620 641.200 ;
      RECT 125.580 1.400 125.860 641.200 ;
      RECT 127.820 1.400 128.100 641.200 ;
      RECT 130.060 1.400 130.340 641.200 ;
      RECT 132.300 1.400 132.580 641.200 ;
      RECT 134.540 1.400 134.820 641.200 ;
      RECT 136.780 1.400 137.060 641.200 ;
      RECT 139.020 1.400 139.300 641.200 ;
      RECT 141.260 1.400 141.540 641.200 ;
      RECT 143.500 1.400 143.780 641.200 ;
      RECT 145.740 1.400 146.020 641.200 ;
      RECT 147.980 1.400 148.260 641.200 ;
      RECT 150.220 1.400 150.500 641.200 ;
      RECT 152.460 1.400 152.740 641.200 ;
      RECT 154.700 1.400 154.980 641.200 ;
      RECT 156.940 1.400 157.220 641.200 ;
      RECT 159.180 1.400 159.460 641.200 ;
      RECT 161.420 1.400 161.700 641.200 ;
      RECT 163.660 1.400 163.940 641.200 ;
      RECT 165.900 1.400 166.180 641.200 ;
      RECT 168.140 1.400 168.420 641.200 ;
      RECT 170.380 1.400 170.660 641.200 ;
      RECT 172.620 1.400 172.900 641.200 ;
      RECT 174.860 1.400 175.140 641.200 ;
      RECT 177.100 1.400 177.380 641.200 ;
      RECT 179.340 1.400 179.620 641.200 ;
      RECT 181.580 1.400 181.860 641.200 ;
      RECT 183.820 1.400 184.100 641.200 ;
      RECT 186.060 1.400 186.340 641.200 ;
      RECT 188.300 1.400 188.580 641.200 ;
      RECT 190.540 1.400 190.820 641.200 ;
      RECT 192.780 1.400 193.060 641.200 ;
      RECT 195.020 1.400 195.300 641.200 ;
      RECT 197.260 1.400 197.540 641.200 ;
      RECT 199.500 1.400 199.780 641.200 ;
      RECT 201.740 1.400 202.020 641.200 ;
      RECT 203.980 1.400 204.260 641.200 ;
      RECT 206.220 1.400 206.500 641.200 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 209.000 642.600 ;
    LAYER metal2 ;
    RECT 0 0 209.000 642.600 ;
    LAYER metal3 ;
    RECT 0.070 0 209.000 642.600 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 7.105 ;
    RECT 0 7.175 0.070 12.845 ;
    RECT 0 12.915 0.070 18.585 ;
    RECT 0 18.655 0.070 24.325 ;
    RECT 0 24.395 0.070 30.065 ;
    RECT 0 30.135 0.070 35.805 ;
    RECT 0 35.875 0.070 41.545 ;
    RECT 0 41.615 0.070 47.285 ;
    RECT 0 47.355 0.070 53.025 ;
    RECT 0 53.095 0.070 58.765 ;
    RECT 0 58.835 0.070 64.505 ;
    RECT 0 64.575 0.070 70.245 ;
    RECT 0 70.315 0.070 75.985 ;
    RECT 0 76.055 0.070 81.725 ;
    RECT 0 81.795 0.070 87.465 ;
    RECT 0 87.535 0.070 93.205 ;
    RECT 0 93.275 0.070 98.945 ;
    RECT 0 99.015 0.070 104.685 ;
    RECT 0 104.755 0.070 110.425 ;
    RECT 0 110.495 0.070 116.165 ;
    RECT 0 116.235 0.070 121.905 ;
    RECT 0 121.975 0.070 127.645 ;
    RECT 0 127.715 0.070 133.385 ;
    RECT 0 133.455 0.070 139.125 ;
    RECT 0 139.195 0.070 144.865 ;
    RECT 0 144.935 0.070 150.605 ;
    RECT 0 150.675 0.070 156.345 ;
    RECT 0 156.415 0.070 162.085 ;
    RECT 0 162.155 0.070 167.825 ;
    RECT 0 167.895 0.070 173.565 ;
    RECT 0 173.635 0.070 179.305 ;
    RECT 0 179.375 0.070 182.805 ;
    RECT 0 182.875 0.070 188.545 ;
    RECT 0 188.615 0.070 194.285 ;
    RECT 0 194.355 0.070 200.025 ;
    RECT 0 200.095 0.070 205.765 ;
    RECT 0 205.835 0.070 211.505 ;
    RECT 0 211.575 0.070 217.245 ;
    RECT 0 217.315 0.070 222.985 ;
    RECT 0 223.055 0.070 228.725 ;
    RECT 0 228.795 0.070 234.465 ;
    RECT 0 234.535 0.070 240.205 ;
    RECT 0 240.275 0.070 245.945 ;
    RECT 0 246.015 0.070 251.685 ;
    RECT 0 251.755 0.070 257.425 ;
    RECT 0 257.495 0.070 263.165 ;
    RECT 0 263.235 0.070 268.905 ;
    RECT 0 268.975 0.070 274.645 ;
    RECT 0 274.715 0.070 280.385 ;
    RECT 0 280.455 0.070 286.125 ;
    RECT 0 286.195 0.070 291.865 ;
    RECT 0 291.935 0.070 297.605 ;
    RECT 0 297.675 0.070 303.345 ;
    RECT 0 303.415 0.070 309.085 ;
    RECT 0 309.155 0.070 314.825 ;
    RECT 0 314.895 0.070 320.565 ;
    RECT 0 320.635 0.070 326.305 ;
    RECT 0 326.375 0.070 332.045 ;
    RECT 0 332.115 0.070 337.785 ;
    RECT 0 337.855 0.070 343.525 ;
    RECT 0 343.595 0.070 349.265 ;
    RECT 0 349.335 0.070 355.005 ;
    RECT 0 355.075 0.070 360.745 ;
    RECT 0 360.815 0.070 364.245 ;
    RECT 0 364.315 0.070 369.985 ;
    RECT 0 370.055 0.070 375.725 ;
    RECT 0 375.795 0.070 381.465 ;
    RECT 0 381.535 0.070 387.205 ;
    RECT 0 387.275 0.070 392.945 ;
    RECT 0 393.015 0.070 398.685 ;
    RECT 0 398.755 0.070 404.425 ;
    RECT 0 404.495 0.070 410.165 ;
    RECT 0 410.235 0.070 415.905 ;
    RECT 0 415.975 0.070 421.645 ;
    RECT 0 421.715 0.070 427.385 ;
    RECT 0 427.455 0.070 433.125 ;
    RECT 0 433.195 0.070 438.865 ;
    RECT 0 438.935 0.070 444.605 ;
    RECT 0 444.675 0.070 450.345 ;
    RECT 0 450.415 0.070 456.085 ;
    RECT 0 456.155 0.070 461.825 ;
    RECT 0 461.895 0.070 467.565 ;
    RECT 0 467.635 0.070 473.305 ;
    RECT 0 473.375 0.070 479.045 ;
    RECT 0 479.115 0.070 484.785 ;
    RECT 0 484.855 0.070 490.525 ;
    RECT 0 490.595 0.070 496.265 ;
    RECT 0 496.335 0.070 502.005 ;
    RECT 0 502.075 0.070 507.745 ;
    RECT 0 507.815 0.070 513.485 ;
    RECT 0 513.555 0.070 519.225 ;
    RECT 0 519.295 0.070 524.965 ;
    RECT 0 525.035 0.070 530.705 ;
    RECT 0 530.775 0.070 536.445 ;
    RECT 0 536.515 0.070 542.185 ;
    RECT 0 542.255 0.070 545.685 ;
    RECT 0 545.755 0.070 551.425 ;
    RECT 0 551.495 0.070 557.165 ;
    RECT 0 557.235 0.070 562.905 ;
    RECT 0 562.975 0.070 568.645 ;
    RECT 0 568.715 0.070 574.385 ;
    RECT 0 574.455 0.070 580.125 ;
    RECT 0 580.195 0.070 585.865 ;
    RECT 0 585.935 0.070 591.605 ;
    RECT 0 591.675 0.070 597.345 ;
    RECT 0 597.415 0.070 600.845 ;
    RECT 0 600.915 0.070 606.585 ;
    RECT 0 606.655 0.070 612.325 ;
    RECT 0 612.395 0.070 642.600 ;
    LAYER metal4 ;
    RECT 0 0 209.000 1.400 ;
    RECT 0 641.200 209.000 642.600 ;
    RECT 0.000 1.400 1.260 641.200 ;
    RECT 1.540 1.400 2.380 641.200 ;
    RECT 2.660 1.400 3.500 641.200 ;
    RECT 3.780 1.400 4.620 641.200 ;
    RECT 4.900 1.400 5.740 641.200 ;
    RECT 6.020 1.400 6.860 641.200 ;
    RECT 7.140 1.400 7.980 641.200 ;
    RECT 8.260 1.400 9.100 641.200 ;
    RECT 9.380 1.400 10.220 641.200 ;
    RECT 10.500 1.400 11.340 641.200 ;
    RECT 11.620 1.400 12.460 641.200 ;
    RECT 12.740 1.400 13.580 641.200 ;
    RECT 13.860 1.400 14.700 641.200 ;
    RECT 14.980 1.400 15.820 641.200 ;
    RECT 16.100 1.400 16.940 641.200 ;
    RECT 17.220 1.400 18.060 641.200 ;
    RECT 18.340 1.400 19.180 641.200 ;
    RECT 19.460 1.400 20.300 641.200 ;
    RECT 20.580 1.400 21.420 641.200 ;
    RECT 21.700 1.400 22.540 641.200 ;
    RECT 22.820 1.400 23.660 641.200 ;
    RECT 23.940 1.400 24.780 641.200 ;
    RECT 25.060 1.400 25.900 641.200 ;
    RECT 26.180 1.400 27.020 641.200 ;
    RECT 27.300 1.400 28.140 641.200 ;
    RECT 28.420 1.400 29.260 641.200 ;
    RECT 29.540 1.400 30.380 641.200 ;
    RECT 30.660 1.400 31.500 641.200 ;
    RECT 31.780 1.400 32.620 641.200 ;
    RECT 32.900 1.400 33.740 641.200 ;
    RECT 34.020 1.400 34.860 641.200 ;
    RECT 35.140 1.400 35.980 641.200 ;
    RECT 36.260 1.400 37.100 641.200 ;
    RECT 37.380 1.400 38.220 641.200 ;
    RECT 38.500 1.400 39.340 641.200 ;
    RECT 39.620 1.400 40.460 641.200 ;
    RECT 40.740 1.400 41.580 641.200 ;
    RECT 41.860 1.400 42.700 641.200 ;
    RECT 42.980 1.400 43.820 641.200 ;
    RECT 44.100 1.400 44.940 641.200 ;
    RECT 45.220 1.400 46.060 641.200 ;
    RECT 46.340 1.400 47.180 641.200 ;
    RECT 47.460 1.400 48.300 641.200 ;
    RECT 48.580 1.400 49.420 641.200 ;
    RECT 49.700 1.400 50.540 641.200 ;
    RECT 50.820 1.400 51.660 641.200 ;
    RECT 51.940 1.400 52.780 641.200 ;
    RECT 53.060 1.400 53.900 641.200 ;
    RECT 54.180 1.400 55.020 641.200 ;
    RECT 55.300 1.400 56.140 641.200 ;
    RECT 56.420 1.400 57.260 641.200 ;
    RECT 57.540 1.400 58.380 641.200 ;
    RECT 58.660 1.400 59.500 641.200 ;
    RECT 59.780 1.400 60.620 641.200 ;
    RECT 60.900 1.400 61.740 641.200 ;
    RECT 62.020 1.400 62.860 641.200 ;
    RECT 63.140 1.400 63.980 641.200 ;
    RECT 64.260 1.400 65.100 641.200 ;
    RECT 65.380 1.400 66.220 641.200 ;
    RECT 66.500 1.400 67.340 641.200 ;
    RECT 67.620 1.400 68.460 641.200 ;
    RECT 68.740 1.400 69.580 641.200 ;
    RECT 69.860 1.400 70.700 641.200 ;
    RECT 70.980 1.400 71.820 641.200 ;
    RECT 72.100 1.400 72.940 641.200 ;
    RECT 73.220 1.400 74.060 641.200 ;
    RECT 74.340 1.400 75.180 641.200 ;
    RECT 75.460 1.400 76.300 641.200 ;
    RECT 76.580 1.400 77.420 641.200 ;
    RECT 77.700 1.400 78.540 641.200 ;
    RECT 78.820 1.400 79.660 641.200 ;
    RECT 79.940 1.400 80.780 641.200 ;
    RECT 81.060 1.400 81.900 641.200 ;
    RECT 82.180 1.400 83.020 641.200 ;
    RECT 83.300 1.400 84.140 641.200 ;
    RECT 84.420 1.400 85.260 641.200 ;
    RECT 85.540 1.400 86.380 641.200 ;
    RECT 86.660 1.400 87.500 641.200 ;
    RECT 87.780 1.400 88.620 641.200 ;
    RECT 88.900 1.400 89.740 641.200 ;
    RECT 90.020 1.400 90.860 641.200 ;
    RECT 91.140 1.400 91.980 641.200 ;
    RECT 92.260 1.400 93.100 641.200 ;
    RECT 93.380 1.400 94.220 641.200 ;
    RECT 94.500 1.400 95.340 641.200 ;
    RECT 95.620 1.400 96.460 641.200 ;
    RECT 96.740 1.400 97.580 641.200 ;
    RECT 97.860 1.400 98.700 641.200 ;
    RECT 98.980 1.400 99.820 641.200 ;
    RECT 100.100 1.400 100.940 641.200 ;
    RECT 101.220 1.400 102.060 641.200 ;
    RECT 102.340 1.400 103.180 641.200 ;
    RECT 103.460 1.400 104.300 641.200 ;
    RECT 104.580 1.400 105.420 641.200 ;
    RECT 105.700 1.400 106.540 641.200 ;
    RECT 106.820 1.400 107.660 641.200 ;
    RECT 107.940 1.400 108.780 641.200 ;
    RECT 109.060 1.400 109.900 641.200 ;
    RECT 110.180 1.400 111.020 641.200 ;
    RECT 111.300 1.400 112.140 641.200 ;
    RECT 112.420 1.400 113.260 641.200 ;
    RECT 113.540 1.400 114.380 641.200 ;
    RECT 114.660 1.400 115.500 641.200 ;
    RECT 115.780 1.400 116.620 641.200 ;
    RECT 116.900 1.400 117.740 641.200 ;
    RECT 118.020 1.400 118.860 641.200 ;
    RECT 119.140 1.400 119.980 641.200 ;
    RECT 120.260 1.400 121.100 641.200 ;
    RECT 121.380 1.400 122.220 641.200 ;
    RECT 122.500 1.400 123.340 641.200 ;
    RECT 123.620 1.400 124.460 641.200 ;
    RECT 124.740 1.400 125.580 641.200 ;
    RECT 125.860 1.400 126.700 641.200 ;
    RECT 126.980 1.400 127.820 641.200 ;
    RECT 128.100 1.400 128.940 641.200 ;
    RECT 129.220 1.400 130.060 641.200 ;
    RECT 130.340 1.400 131.180 641.200 ;
    RECT 131.460 1.400 132.300 641.200 ;
    RECT 132.580 1.400 133.420 641.200 ;
    RECT 133.700 1.400 134.540 641.200 ;
    RECT 134.820 1.400 135.660 641.200 ;
    RECT 135.940 1.400 136.780 641.200 ;
    RECT 137.060 1.400 137.900 641.200 ;
    RECT 138.180 1.400 139.020 641.200 ;
    RECT 139.300 1.400 140.140 641.200 ;
    RECT 140.420 1.400 141.260 641.200 ;
    RECT 141.540 1.400 142.380 641.200 ;
    RECT 142.660 1.400 143.500 641.200 ;
    RECT 143.780 1.400 144.620 641.200 ;
    RECT 144.900 1.400 145.740 641.200 ;
    RECT 146.020 1.400 146.860 641.200 ;
    RECT 147.140 1.400 147.980 641.200 ;
    RECT 148.260 1.400 149.100 641.200 ;
    RECT 149.380 1.400 150.220 641.200 ;
    RECT 150.500 1.400 151.340 641.200 ;
    RECT 151.620 1.400 152.460 641.200 ;
    RECT 152.740 1.400 153.580 641.200 ;
    RECT 153.860 1.400 154.700 641.200 ;
    RECT 154.980 1.400 155.820 641.200 ;
    RECT 156.100 1.400 156.940 641.200 ;
    RECT 157.220 1.400 158.060 641.200 ;
    RECT 158.340 1.400 159.180 641.200 ;
    RECT 159.460 1.400 160.300 641.200 ;
    RECT 160.580 1.400 161.420 641.200 ;
    RECT 161.700 1.400 162.540 641.200 ;
    RECT 162.820 1.400 163.660 641.200 ;
    RECT 163.940 1.400 164.780 641.200 ;
    RECT 165.060 1.400 165.900 641.200 ;
    RECT 166.180 1.400 167.020 641.200 ;
    RECT 167.300 1.400 168.140 641.200 ;
    RECT 168.420 1.400 169.260 641.200 ;
    RECT 169.540 1.400 170.380 641.200 ;
    RECT 170.660 1.400 171.500 641.200 ;
    RECT 171.780 1.400 172.620 641.200 ;
    RECT 172.900 1.400 173.740 641.200 ;
    RECT 174.020 1.400 174.860 641.200 ;
    RECT 175.140 1.400 175.980 641.200 ;
    RECT 176.260 1.400 177.100 641.200 ;
    RECT 177.380 1.400 178.220 641.200 ;
    RECT 178.500 1.400 179.340 641.200 ;
    RECT 179.620 1.400 180.460 641.200 ;
    RECT 180.740 1.400 181.580 641.200 ;
    RECT 181.860 1.400 182.700 641.200 ;
    RECT 182.980 1.400 183.820 641.200 ;
    RECT 184.100 1.400 184.940 641.200 ;
    RECT 185.220 1.400 186.060 641.200 ;
    RECT 186.340 1.400 187.180 641.200 ;
    RECT 187.460 1.400 188.300 641.200 ;
    RECT 188.580 1.400 189.420 641.200 ;
    RECT 189.700 1.400 190.540 641.200 ;
    RECT 190.820 1.400 191.660 641.200 ;
    RECT 191.940 1.400 192.780 641.200 ;
    RECT 193.060 1.400 193.900 641.200 ;
    RECT 194.180 1.400 195.020 641.200 ;
    RECT 195.300 1.400 196.140 641.200 ;
    RECT 196.420 1.400 197.260 641.200 ;
    RECT 197.540 1.400 198.380 641.200 ;
    RECT 198.660 1.400 199.500 641.200 ;
    RECT 199.780 1.400 200.620 641.200 ;
    RECT 200.900 1.400 201.740 641.200 ;
    RECT 202.020 1.400 202.860 641.200 ;
    RECT 203.140 1.400 203.980 641.200 ;
    RECT 204.260 1.400 205.100 641.200 ;
    RECT 205.380 1.400 206.220 641.200 ;
    RECT 206.500 1.400 207.340 641.200 ;
    RECT 207.620 1.400 209.000 641.200 ;
    LAYER OVERLAP ;
    RECT 0 0 209.000 642.600 ;
  END
END sram_32x1024_2r1w

END LIBRARY
