VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_32x128_2r1w
  FOREIGN fakeram_32x128_2r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 16.589 BY 10.368 ;
  CLASS BLOCK ;
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.276 0.024 0.300 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.756 0.024 0.780 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.236 0.024 1.260 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.716 0.024 1.740 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.196 0.024 2.220 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.676 0.024 2.700 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.156 0.024 3.180 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.636 0.024 3.660 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 0.276 16.589 0.300 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 0.756 16.589 0.780 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 1.236 16.589 1.260 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 1.716 16.589 1.740 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 2.196 16.589 2.220 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 2.676 16.589 2.700 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 3.156 16.589 3.180 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 3.636 16.589 3.660 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 0.000 0.225 0.018 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.531 0.000 0.549 0.018 ;
    END
  END w0_wd_in[17]
  PIN w0_wd_in[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.855 0.000 0.873 0.018 ;
    END
  END w0_wd_in[18]
  PIN w0_wd_in[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.179 0.000 1.197 0.018 ;
    END
  END w0_wd_in[19]
  PIN w0_wd_in[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.503 0.000 1.521 0.018 ;
    END
  END w0_wd_in[20]
  PIN w0_wd_in[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.827 0.000 1.845 0.018 ;
    END
  END w0_wd_in[21]
  PIN w0_wd_in[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.151 0.000 2.169 0.018 ;
    END
  END w0_wd_in[22]
  PIN w0_wd_in[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.475 0.000 2.493 0.018 ;
    END
  END w0_wd_in[23]
  PIN w0_wd_in[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.799 0.000 2.817 0.018 ;
    END
  END w0_wd_in[24]
  PIN w0_wd_in[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.123 0.000 3.141 0.018 ;
    END
  END w0_wd_in[25]
  PIN w0_wd_in[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.447 0.000 3.465 0.018 ;
    END
  END w0_wd_in[26]
  PIN w0_wd_in[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.771 0.000 3.789 0.018 ;
    END
  END w0_wd_in[27]
  PIN w0_wd_in[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.095 0.000 4.113 0.018 ;
    END
  END w0_wd_in[28]
  PIN w0_wd_in[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.419 0.000 4.437 0.018 ;
    END
  END w0_wd_in[29]
  PIN w0_wd_in[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.743 0.000 4.761 0.018 ;
    END
  END w0_wd_in[30]
  PIN w0_wd_in[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.067 0.000 5.085 0.018 ;
    END
  END w0_wd_in[31]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.391 0.000 5.409 0.018 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.715 0.000 5.733 0.018 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.039 0.000 6.057 0.018 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.363 0.000 6.381 0.018 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.687 0.000 6.705 0.018 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.011 0.000 7.029 0.018 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.335 0.000 7.353 0.018 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.659 0.000 7.677 0.018 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.983 0.000 8.001 0.018 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.307 0.000 8.325 0.018 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.631 0.000 8.649 0.018 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.955 0.000 8.973 0.018 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.279 0.000 9.297 0.018 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.603 0.000 9.621 0.018 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.927 0.000 9.945 0.018 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.251 0.000 10.269 0.018 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 10.350 0.225 10.368 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.603 10.350 0.621 10.368 ;
    END
  END r0_rd_out[17]
  PIN r0_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.999 10.350 1.017 10.368 ;
    END
  END r0_rd_out[18]
  PIN r0_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.395 10.350 1.413 10.368 ;
    END
  END r0_rd_out[19]
  PIN r0_rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.791 10.350 1.809 10.368 ;
    END
  END r0_rd_out[20]
  PIN r0_rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.187 10.350 2.205 10.368 ;
    END
  END r0_rd_out[21]
  PIN r0_rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.583 10.350 2.601 10.368 ;
    END
  END r0_rd_out[22]
  PIN r0_rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.979 10.350 2.997 10.368 ;
    END
  END r0_rd_out[23]
  PIN r0_rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.375 10.350 3.393 10.368 ;
    END
  END r0_rd_out[24]
  PIN r0_rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.771 10.350 3.789 10.368 ;
    END
  END r0_rd_out[25]
  PIN r0_rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.167 10.350 4.185 10.368 ;
    END
  END r0_rd_out[26]
  PIN r0_rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.563 10.350 4.581 10.368 ;
    END
  END r0_rd_out[27]
  PIN r0_rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.959 10.350 4.977 10.368 ;
    END
  END r0_rd_out[28]
  PIN r0_rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.355 10.350 5.373 10.368 ;
    END
  END r0_rd_out[29]
  PIN r0_rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.751 10.350 5.769 10.368 ;
    END
  END r0_rd_out[30]
  PIN r0_rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.147 10.350 6.165 10.368 ;
    END
  END r0_rd_out[31]
  PIN r1_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.575 0.000 10.593 0.018 ;
    END
  END r1_rd_out[0]
  PIN r1_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.899 0.000 10.917 0.018 ;
    END
  END r1_rd_out[1]
  PIN r1_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 11.223 0.000 11.241 0.018 ;
    END
  END r1_rd_out[2]
  PIN r1_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 11.547 0.000 11.565 0.018 ;
    END
  END r1_rd_out[3]
  PIN r1_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 11.871 0.000 11.889 0.018 ;
    END
  END r1_rd_out[4]
  PIN r1_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.195 0.000 12.213 0.018 ;
    END
  END r1_rd_out[5]
  PIN r1_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.519 0.000 12.537 0.018 ;
    END
  END r1_rd_out[6]
  PIN r1_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.843 0.000 12.861 0.018 ;
    END
  END r1_rd_out[7]
  PIN r1_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 13.167 0.000 13.185 0.018 ;
    END
  END r1_rd_out[8]
  PIN r1_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 13.491 0.000 13.509 0.018 ;
    END
  END r1_rd_out[9]
  PIN r1_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 13.815 0.000 13.833 0.018 ;
    END
  END r1_rd_out[10]
  PIN r1_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 14.139 0.000 14.157 0.018 ;
    END
  END r1_rd_out[11]
  PIN r1_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 14.463 0.000 14.481 0.018 ;
    END
  END r1_rd_out[12]
  PIN r1_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 14.787 0.000 14.805 0.018 ;
    END
  END r1_rd_out[13]
  PIN r1_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 15.111 0.000 15.129 0.018 ;
    END
  END r1_rd_out[14]
  PIN r1_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 15.435 0.000 15.453 0.018 ;
    END
  END r1_rd_out[15]
  PIN r1_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.543 10.350 6.561 10.368 ;
    END
  END r1_rd_out[16]
  PIN r1_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.939 10.350 6.957 10.368 ;
    END
  END r1_rd_out[17]
  PIN r1_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.335 10.350 7.353 10.368 ;
    END
  END r1_rd_out[18]
  PIN r1_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.731 10.350 7.749 10.368 ;
    END
  END r1_rd_out[19]
  PIN r1_rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.127 10.350 8.145 10.368 ;
    END
  END r1_rd_out[20]
  PIN r1_rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.523 10.350 8.541 10.368 ;
    END
  END r1_rd_out[21]
  PIN r1_rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.919 10.350 8.937 10.368 ;
    END
  END r1_rd_out[22]
  PIN r1_rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.315 10.350 9.333 10.368 ;
    END
  END r1_rd_out[23]
  PIN r1_rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.711 10.350 9.729 10.368 ;
    END
  END r1_rd_out[24]
  PIN r1_rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.107 10.350 10.125 10.368 ;
    END
  END r1_rd_out[25]
  PIN r1_rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.503 10.350 10.521 10.368 ;
    END
  END r1_rd_out[26]
  PIN r1_rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.899 10.350 10.917 10.368 ;
    END
  END r1_rd_out[27]
  PIN r1_rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 11.295 10.350 11.313 10.368 ;
    END
  END r1_rd_out[28]
  PIN r1_rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 11.691 10.350 11.709 10.368 ;
    END
  END r1_rd_out[29]
  PIN r1_rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.087 10.350 12.105 10.368 ;
    END
  END r1_rd_out[30]
  PIN r1_rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.483 10.350 12.501 10.368 ;
    END
  END r1_rd_out[31]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.116 0.024 4.140 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.596 0.024 4.620 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.076 0.024 5.100 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.556 0.024 5.580 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 4.116 16.589 4.140 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 4.596 16.589 4.620 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 5.076 16.589 5.100 ;
    END
  END w0_addr_in[6]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.036 0.024 6.060 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.516 0.024 6.540 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.996 0.024 7.020 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.476 0.024 7.500 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 5.556 16.589 5.580 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 6.036 16.589 6.060 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 6.516 16.589 6.540 ;
    END
  END r0_addr_in[6]
  PIN r1_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.956 0.024 7.980 ;
    END
  END r1_addr_in[0]
  PIN r1_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.436 0.024 8.460 ;
    END
  END r1_addr_in[1]
  PIN r1_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.916 0.024 8.940 ;
    END
  END r1_addr_in[2]
  PIN r1_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.396 0.024 9.420 ;
    END
  END r1_addr_in[3]
  PIN r1_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 6.996 16.589 7.020 ;
    END
  END r1_addr_in[4]
  PIN r1_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 7.476 16.589 7.500 ;
    END
  END r1_addr_in[5]
  PIN r1_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.565 7.956 16.589 7.980 ;
    END
  END r1_addr_in[6]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.879 10.350 12.897 10.368 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 13.275 10.350 13.293 10.368 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 13.671 10.350 13.689 10.368 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 14.067 10.350 14.085 10.368 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 14.463 10.350 14.481 10.368 ;
    END
  END r0_clk
  PIN r1_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 14.859 10.350 14.877 10.368 ;
    END
  END r1_ce_in
  PIN r1_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 15.255 10.350 15.273 10.368 ;
    END
  END r1_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.108 0.192 16.481 0.288 ;
      RECT 0.108 0.960 16.481 1.056 ;
      RECT 0.108 1.728 16.481 1.824 ;
      RECT 0.108 2.496 16.481 2.592 ;
      RECT 0.108 3.264 16.481 3.360 ;
      RECT 0.108 4.032 16.481 4.128 ;
      RECT 0.108 4.800 16.481 4.896 ;
      RECT 0.108 5.568 16.481 5.664 ;
      RECT 0.108 6.336 16.481 6.432 ;
      RECT 0.108 7.104 16.481 7.200 ;
      RECT 0.108 7.872 16.481 7.968 ;
      RECT 0.108 8.640 16.481 8.736 ;
      RECT 0.108 9.408 16.481 9.504 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.108 0.192 16.481 0.288 ;
      RECT 0.108 0.960 16.481 1.056 ;
      RECT 0.108 1.728 16.481 1.824 ;
      RECT 0.108 2.496 16.481 2.592 ;
      RECT 0.108 3.264 16.481 3.360 ;
      RECT 0.108 4.032 16.481 4.128 ;
      RECT 0.108 4.800 16.481 4.896 ;
      RECT 0.108 5.568 16.481 5.664 ;
      RECT 0.108 6.336 16.481 6.432 ;
      RECT 0.108 7.104 16.481 7.200 ;
      RECT 0.108 7.872 16.481 7.968 ;
      RECT 0.108 8.640 16.481 8.736 ;
      RECT 0.108 9.408 16.481 9.504 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 16.589 10.368 ;
    LAYER M2 ;
    RECT 0 0 16.589 10.368 ;
    LAYER M3 ;
    RECT 0 0 16.589 10.368 ;
    LAYER M4 ;
    RECT 0 0 16.589 10.368 ;
  END
END fakeram_32x128_2r1w

END LIBRARY
