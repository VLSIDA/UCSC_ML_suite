VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_18x256_1r1w
  FOREIGN fakeram_18x256_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 388.240 BY 323.680 ;
  CLASS BLOCK ;
  PIN w0_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 6.650 0.800 6.950 ;
    END
  END w0_mask_in[0]
  PIN w0_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.810 0.800 15.110 ;
    END
  END w0_mask_in[1]
  PIN w0_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.970 0.800 23.270 ;
    END
  END w0_mask_in[2]
  PIN w0_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.130 0.800 31.430 ;
    END
  END w0_mask_in[3]
  PIN w0_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.290 0.800 39.590 ;
    END
  END w0_mask_in[4]
  PIN w0_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 47.450 0.800 47.750 ;
    END
  END w0_mask_in[5]
  PIN w0_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.610 0.800 55.910 ;
    END
  END w0_mask_in[6]
  PIN w0_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 63.770 0.800 64.070 ;
    END
  END w0_mask_in[7]
  PIN w0_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.930 0.800 72.230 ;
    END
  END w0_mask_in[8]
  PIN w0_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 80.090 0.800 80.390 ;
    END
  END w0_mask_in[9]
  PIN w0_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 88.250 0.800 88.550 ;
    END
  END w0_mask_in[10]
  PIN w0_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 96.410 0.800 96.710 ;
    END
  END w0_mask_in[11]
  PIN w0_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 104.570 0.800 104.870 ;
    END
  END w0_mask_in[12]
  PIN w0_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 112.730 0.800 113.030 ;
    END
  END w0_mask_in[13]
  PIN w0_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 120.890 0.800 121.190 ;
    END
  END w0_mask_in[14]
  PIN w0_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 129.050 0.800 129.350 ;
    END
  END w0_mask_in[15]
  PIN w0_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 137.210 0.800 137.510 ;
    END
  END w0_mask_in[16]
  PIN w0_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 145.370 0.800 145.670 ;
    END
  END w0_mask_in[17]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 152.850 0.800 153.150 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 161.010 0.800 161.310 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 169.170 0.800 169.470 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 177.330 0.800 177.630 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 185.490 0.800 185.790 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 193.650 0.800 193.950 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 201.810 0.800 202.110 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 209.970 0.800 210.270 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 218.130 0.800 218.430 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 226.290 0.800 226.590 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 234.450 0.800 234.750 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 242.610 0.800 242.910 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 250.770 0.800 251.070 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 258.930 0.800 259.230 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 267.090 0.800 267.390 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 275.250 0.800 275.550 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 283.410 0.800 283.710 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 291.570 0.800 291.870 ;
    END
  END w0_wd_in[17]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 0.000 4.670 0.350 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 25.230 0.000 25.370 0.350 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 45.930 0.000 46.070 0.350 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 66.630 0.000 66.770 0.350 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 87.330 0.000 87.470 0.350 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 108.030 0.000 108.170 0.350 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 128.730 0.000 128.870 0.350 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 149.430 0.000 149.570 0.350 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 170.130 0.000 170.270 0.350 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 190.830 0.000 190.970 0.350 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 211.530 0.000 211.670 0.350 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 232.230 0.000 232.370 0.350 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 252.930 0.000 253.070 0.350 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 273.630 0.000 273.770 0.350 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 294.330 0.000 294.470 0.350 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 315.030 0.000 315.170 0.350 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 335.730 0.000 335.870 0.350 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 356.430 0.000 356.570 0.350 ;
    END
  END r0_rd_out[17]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 387.440 6.650 388.240 6.950 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 387.440 20.930 388.240 21.230 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 387.440 35.210 388.240 35.510 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 387.440 49.490 388.240 49.790 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 387.440 63.770 388.240 64.070 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 387.440 78.050 388.240 78.350 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 387.440 92.330 388.240 92.630 ;
    END
  END w0_addr_in[6]
  PIN w0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 387.440 106.610 388.240 106.910 ;
    END
  END w0_addr_in[7]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 323.330 4.670 323.680 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 23.390 323.330 23.530 323.680 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 42.250 323.330 42.390 323.680 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 61.110 323.330 61.250 323.680 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 79.970 323.330 80.110 323.680 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 98.830 323.330 98.970 323.680 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 117.690 323.330 117.830 323.680 ;
    END
  END r0_addr_in[6]
  PIN r0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 136.550 323.330 136.690 323.680 ;
    END
  END r0_addr_in[7]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 387.440 111.370 388.240 111.670 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 387.440 116.130 388.240 116.430 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 387.440 120.890 388.240 121.190 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 137.470 323.330 137.610 323.680 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 138.390 323.330 138.530 323.680 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 3.240 6.800 5.960 316.880 ;
      RECT 14.120 6.800 16.840 316.880 ;
      RECT 25.000 6.800 27.720 316.880 ;
      RECT 35.880 6.800 38.600 316.880 ;
      RECT 46.760 6.800 49.480 316.880 ;
      RECT 57.640 6.800 60.360 316.880 ;
      RECT 68.520 6.800 71.240 316.880 ;
      RECT 79.400 6.800 82.120 316.880 ;
      RECT 90.280 6.800 93.000 316.880 ;
      RECT 101.160 6.800 103.880 316.880 ;
      RECT 112.040 6.800 114.760 316.880 ;
      RECT 122.920 6.800 125.640 316.880 ;
      RECT 133.800 6.800 136.520 316.880 ;
      RECT 144.680 6.800 147.400 316.880 ;
      RECT 155.560 6.800 158.280 316.880 ;
      RECT 166.440 6.800 169.160 316.880 ;
      RECT 177.320 6.800 180.040 316.880 ;
      RECT 188.200 6.800 190.920 316.880 ;
      RECT 199.080 6.800 201.800 316.880 ;
      RECT 209.960 6.800 212.680 316.880 ;
      RECT 220.840 6.800 223.560 316.880 ;
      RECT 231.720 6.800 234.440 316.880 ;
      RECT 242.600 6.800 245.320 316.880 ;
      RECT 253.480 6.800 256.200 316.880 ;
      RECT 264.360 6.800 267.080 316.880 ;
      RECT 275.240 6.800 277.960 316.880 ;
      RECT 286.120 6.800 288.840 316.880 ;
      RECT 297.000 6.800 299.720 316.880 ;
      RECT 307.880 6.800 310.600 316.880 ;
      RECT 318.760 6.800 321.480 316.880 ;
      RECT 329.640 6.800 332.360 316.880 ;
      RECT 340.520 6.800 343.240 316.880 ;
      RECT 351.400 6.800 354.120 316.880 ;
      RECT 362.280 6.800 365.000 316.880 ;
      RECT 373.160 6.800 375.880 316.880 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 8.680 6.800 11.400 316.880 ;
      RECT 19.560 6.800 22.280 316.880 ;
      RECT 30.440 6.800 33.160 316.880 ;
      RECT 41.320 6.800 44.040 316.880 ;
      RECT 52.200 6.800 54.920 316.880 ;
      RECT 63.080 6.800 65.800 316.880 ;
      RECT 73.960 6.800 76.680 316.880 ;
      RECT 84.840 6.800 87.560 316.880 ;
      RECT 95.720 6.800 98.440 316.880 ;
      RECT 106.600 6.800 109.320 316.880 ;
      RECT 117.480 6.800 120.200 316.880 ;
      RECT 128.360 6.800 131.080 316.880 ;
      RECT 139.240 6.800 141.960 316.880 ;
      RECT 150.120 6.800 152.840 316.880 ;
      RECT 161.000 6.800 163.720 316.880 ;
      RECT 171.880 6.800 174.600 316.880 ;
      RECT 182.760 6.800 185.480 316.880 ;
      RECT 193.640 6.800 196.360 316.880 ;
      RECT 204.520 6.800 207.240 316.880 ;
      RECT 215.400 6.800 218.120 316.880 ;
      RECT 226.280 6.800 229.000 316.880 ;
      RECT 237.160 6.800 239.880 316.880 ;
      RECT 248.040 6.800 250.760 316.880 ;
      RECT 258.920 6.800 261.640 316.880 ;
      RECT 269.800 6.800 272.520 316.880 ;
      RECT 280.680 6.800 283.400 316.880 ;
      RECT 291.560 6.800 294.280 316.880 ;
      RECT 302.440 6.800 305.160 316.880 ;
      RECT 313.320 6.800 316.040 316.880 ;
      RECT 324.200 6.800 326.920 316.880 ;
      RECT 335.080 6.800 337.800 316.880 ;
      RECT 345.960 6.800 348.680 316.880 ;
      RECT 356.840 6.800 359.560 316.880 ;
      RECT 367.720 6.800 370.440 316.880 ;
      RECT 378.600 6.800 381.320 316.880 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 388.240 323.680 ;
    LAYER met2 ;
    RECT 0 0 388.240 323.680 ;
    LAYER met3 ;
    RECT 0.800 0 388.240 323.680 ;
    LAYER met4 ;
    RECT 0 0 388.240 6.800 ;
    RECT 0 316.880 388.240 323.680 ;
    RECT 0.000 6.800 3.240 316.880 ;
    RECT 5.960 6.800 8.680 316.880 ;
    RECT 11.400 6.800 14.120 316.880 ;
    RECT 16.840 6.800 19.560 316.880 ;
    RECT 22.280 6.800 25.000 316.880 ;
    RECT 27.720 6.800 30.440 316.880 ;
    RECT 33.160 6.800 35.880 316.880 ;
    RECT 38.600 6.800 41.320 316.880 ;
    RECT 44.040 6.800 46.760 316.880 ;
    RECT 49.480 6.800 52.200 316.880 ;
    RECT 54.920 6.800 57.640 316.880 ;
    RECT 60.360 6.800 63.080 316.880 ;
    RECT 65.800 6.800 68.520 316.880 ;
    RECT 71.240 6.800 73.960 316.880 ;
    RECT 76.680 6.800 79.400 316.880 ;
    RECT 82.120 6.800 84.840 316.880 ;
    RECT 87.560 6.800 90.280 316.880 ;
    RECT 93.000 6.800 95.720 316.880 ;
    RECT 98.440 6.800 101.160 316.880 ;
    RECT 103.880 6.800 106.600 316.880 ;
    RECT 109.320 6.800 112.040 316.880 ;
    RECT 114.760 6.800 117.480 316.880 ;
    RECT 120.200 6.800 122.920 316.880 ;
    RECT 125.640 6.800 128.360 316.880 ;
    RECT 131.080 6.800 133.800 316.880 ;
    RECT 136.520 6.800 139.240 316.880 ;
    RECT 141.960 6.800 144.680 316.880 ;
    RECT 147.400 6.800 150.120 316.880 ;
    RECT 152.840 6.800 155.560 316.880 ;
    RECT 158.280 6.800 161.000 316.880 ;
    RECT 163.720 6.800 166.440 316.880 ;
    RECT 169.160 6.800 171.880 316.880 ;
    RECT 174.600 6.800 177.320 316.880 ;
    RECT 180.040 6.800 182.760 316.880 ;
    RECT 185.480 6.800 188.200 316.880 ;
    RECT 190.920 6.800 193.640 316.880 ;
    RECT 196.360 6.800 199.080 316.880 ;
    RECT 201.800 6.800 204.520 316.880 ;
    RECT 207.240 6.800 209.960 316.880 ;
    RECT 212.680 6.800 215.400 316.880 ;
    RECT 218.120 6.800 220.840 316.880 ;
    RECT 223.560 6.800 226.280 316.880 ;
    RECT 229.000 6.800 231.720 316.880 ;
    RECT 234.440 6.800 237.160 316.880 ;
    RECT 239.880 6.800 242.600 316.880 ;
    RECT 245.320 6.800 248.040 316.880 ;
    RECT 250.760 6.800 253.480 316.880 ;
    RECT 256.200 6.800 258.920 316.880 ;
    RECT 261.640 6.800 264.360 316.880 ;
    RECT 267.080 6.800 269.800 316.880 ;
    RECT 272.520 6.800 275.240 316.880 ;
    RECT 277.960 6.800 280.680 316.880 ;
    RECT 283.400 6.800 286.120 316.880 ;
    RECT 288.840 6.800 291.560 316.880 ;
    RECT 294.280 6.800 297.000 316.880 ;
    RECT 299.720 6.800 302.440 316.880 ;
    RECT 305.160 6.800 307.880 316.880 ;
    RECT 310.600 6.800 313.320 316.880 ;
    RECT 316.040 6.800 318.760 316.880 ;
    RECT 321.480 6.800 324.200 316.880 ;
    RECT 326.920 6.800 329.640 316.880 ;
    RECT 332.360 6.800 335.080 316.880 ;
    RECT 337.800 6.800 340.520 316.880 ;
    RECT 343.240 6.800 345.960 316.880 ;
    RECT 348.680 6.800 351.400 316.880 ;
    RECT 354.120 6.800 356.840 316.880 ;
    RECT 359.560 6.800 362.280 316.880 ;
    RECT 365.000 6.800 367.720 316.880 ;
    RECT 370.440 6.800 373.160 316.880 ;
    RECT 375.880 6.800 378.600 316.880 ;
    RECT 381.320 6.800 388.240 316.880 ;
    LAYER OVERLAP ;
    RECT 0 0 388.240 323.680 ;
  END
END fakeram_18x256_1r1w

END LIBRARY
