VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_1x256_1r1w
  FOREIGN fakeram_1x256_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 229.540 BY 484.160 ;
  CLASS BLOCK ;
  PIN w0_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 6.650 0.800 6.950 ;
    END
  END w0_mask_in[0]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 7.330 0.800 7.630 ;
    END
  END w0_wd_in[0]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 0.000 4.670 0.350 ;
    END
  END r0_rd_out[0]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 228.740 6.650 229.540 6.950 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 228.740 123.610 229.540 123.910 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 228.740 240.570 229.540 240.870 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 228.740 357.530 229.540 357.830 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 228.740 474.490 229.540 474.790 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 228.740 591.450 229.540 591.750 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 228.740 708.410 229.540 708.710 ;
    END
  END w0_addr_in[6]
  PIN w0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 228.740 825.370 229.540 825.670 ;
    END
  END w0_addr_in[7]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 483.810 4.670 484.160 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 77.670 483.810 77.810 484.160 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 150.810 483.810 150.950 484.160 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 223.950 483.810 224.090 484.160 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 297.090 483.810 297.230 484.160 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 370.230 483.810 370.370 484.160 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 443.370 483.810 443.510 484.160 ;
    END
  END r0_addr_in[6]
  PIN r0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 516.510 483.810 516.650 484.160 ;
    END
  END r0_addr_in[7]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 228.740 826.730 229.540 827.030 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 228.740 828.090 229.540 828.390 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 228.740 829.450 229.540 829.750 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 516.970 483.810 517.110 484.160 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 517.430 483.810 517.570 484.160 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 3.240 6.800 5.960 477.360 ;
      RECT 14.120 6.800 16.840 477.360 ;
      RECT 25.000 6.800 27.720 477.360 ;
      RECT 35.880 6.800 38.600 477.360 ;
      RECT 46.760 6.800 49.480 477.360 ;
      RECT 57.640 6.800 60.360 477.360 ;
      RECT 68.520 6.800 71.240 477.360 ;
      RECT 79.400 6.800 82.120 477.360 ;
      RECT 90.280 6.800 93.000 477.360 ;
      RECT 101.160 6.800 103.880 477.360 ;
      RECT 112.040 6.800 114.760 477.360 ;
      RECT 122.920 6.800 125.640 477.360 ;
      RECT 133.800 6.800 136.520 477.360 ;
      RECT 144.680 6.800 147.400 477.360 ;
      RECT 155.560 6.800 158.280 477.360 ;
      RECT 166.440 6.800 169.160 477.360 ;
      RECT 177.320 6.800 180.040 477.360 ;
      RECT 188.200 6.800 190.920 477.360 ;
      RECT 199.080 6.800 201.800 477.360 ;
      RECT 209.960 6.800 212.680 477.360 ;
      RECT 220.840 6.800 223.560 477.360 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 8.680 6.800 11.400 477.360 ;
      RECT 19.560 6.800 22.280 477.360 ;
      RECT 30.440 6.800 33.160 477.360 ;
      RECT 41.320 6.800 44.040 477.360 ;
      RECT 52.200 6.800 54.920 477.360 ;
      RECT 63.080 6.800 65.800 477.360 ;
      RECT 73.960 6.800 76.680 477.360 ;
      RECT 84.840 6.800 87.560 477.360 ;
      RECT 95.720 6.800 98.440 477.360 ;
      RECT 106.600 6.800 109.320 477.360 ;
      RECT 117.480 6.800 120.200 477.360 ;
      RECT 128.360 6.800 131.080 477.360 ;
      RECT 139.240 6.800 141.960 477.360 ;
      RECT 150.120 6.800 152.840 477.360 ;
      RECT 161.000 6.800 163.720 477.360 ;
      RECT 171.880 6.800 174.600 477.360 ;
      RECT 182.760 6.800 185.480 477.360 ;
      RECT 193.640 6.800 196.360 477.360 ;
      RECT 204.520 6.800 207.240 477.360 ;
      RECT 215.400 6.800 218.120 477.360 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 229.540 484.160 ;
    LAYER met2 ;
    RECT 0 0 229.540 484.160 ;
    LAYER met3 ;
    RECT 0.800 0 229.540 484.160 ;
    LAYER met4 ;
    RECT 0 0 229.540 6.800 ;
    RECT 0 477.360 229.540 484.160 ;
    RECT 0.000 6.800 3.240 477.360 ;
    RECT 5.960 6.800 8.680 477.360 ;
    RECT 11.400 6.800 14.120 477.360 ;
    RECT 16.840 6.800 19.560 477.360 ;
    RECT 22.280 6.800 25.000 477.360 ;
    RECT 27.720 6.800 30.440 477.360 ;
    RECT 33.160 6.800 35.880 477.360 ;
    RECT 38.600 6.800 41.320 477.360 ;
    RECT 44.040 6.800 46.760 477.360 ;
    RECT 49.480 6.800 52.200 477.360 ;
    RECT 54.920 6.800 57.640 477.360 ;
    RECT 60.360 6.800 63.080 477.360 ;
    RECT 65.800 6.800 68.520 477.360 ;
    RECT 71.240 6.800 73.960 477.360 ;
    RECT 76.680 6.800 79.400 477.360 ;
    RECT 82.120 6.800 84.840 477.360 ;
    RECT 87.560 6.800 90.280 477.360 ;
    RECT 93.000 6.800 95.720 477.360 ;
    RECT 98.440 6.800 101.160 477.360 ;
    RECT 103.880 6.800 106.600 477.360 ;
    RECT 109.320 6.800 112.040 477.360 ;
    RECT 114.760 6.800 117.480 477.360 ;
    RECT 120.200 6.800 122.920 477.360 ;
    RECT 125.640 6.800 128.360 477.360 ;
    RECT 131.080 6.800 133.800 477.360 ;
    RECT 136.520 6.800 139.240 477.360 ;
    RECT 141.960 6.800 144.680 477.360 ;
    RECT 147.400 6.800 150.120 477.360 ;
    RECT 152.840 6.800 155.560 477.360 ;
    RECT 158.280 6.800 161.000 477.360 ;
    RECT 163.720 6.800 166.440 477.360 ;
    RECT 169.160 6.800 171.880 477.360 ;
    RECT 174.600 6.800 177.320 477.360 ;
    RECT 180.040 6.800 182.760 477.360 ;
    RECT 185.480 6.800 188.200 477.360 ;
    RECT 190.920 6.800 193.640 477.360 ;
    RECT 196.360 6.800 199.080 477.360 ;
    RECT 201.800 6.800 204.520 477.360 ;
    RECT 207.240 6.800 209.960 477.360 ;
    RECT 212.680 6.800 215.400 477.360 ;
    RECT 218.120 6.800 220.840 477.360 ;
    RECT 223.560 6.800 229.540 477.360 ;
    LAYER OVERLAP ;
    RECT 0 0 229.540 484.160 ;
  END
END fakeram_1x256_1r1w

END LIBRARY
