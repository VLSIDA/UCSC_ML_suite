VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_32x1024_1r1w
  FOREIGN sram_32x1024_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 159.980 BY 485.800 ;
  CLASS BLOCK ;
  PIN w_mask_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 -0.595 0.070 -0.525 ;
    END
  END w_mask_w1[0]
  PIN w_mask_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_w1[1]
  PIN w_mask_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_w1[2]
  PIN w_mask_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.425 0.070 12.495 ;
    END
  END w_mask_w1[3]
  PIN w_mask_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_w1[4]
  PIN w_mask_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.105 0.070 21.175 ;
    END
  END w_mask_w1[5]
  PIN w_mask_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.445 0.070 25.515 ;
    END
  END w_mask_w1[6]
  PIN w_mask_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END w_mask_w1[7]
  PIN w_mask_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.125 0.070 34.195 ;
    END
  END w_mask_w1[8]
  PIN w_mask_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.465 0.070 38.535 ;
    END
  END w_mask_w1[9]
  PIN w_mask_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END w_mask_w1[10]
  PIN w_mask_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.145 0.070 47.215 ;
    END
  END w_mask_w1[11]
  PIN w_mask_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.485 0.070 51.555 ;
    END
  END w_mask_w1[12]
  PIN w_mask_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END w_mask_w1[13]
  PIN w_mask_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_w1[14]
  PIN w_mask_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.505 0.070 64.575 ;
    END
  END w_mask_w1[15]
  PIN w_mask_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END w_mask_w1[16]
  PIN w_mask_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.185 0.070 73.255 ;
    END
  END w_mask_w1[17]
  PIN w_mask_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.525 0.070 77.595 ;
    END
  END w_mask_w1[18]
  PIN w_mask_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END w_mask_w1[19]
  PIN w_mask_w1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.205 0.070 86.275 ;
    END
  END w_mask_w1[20]
  PIN w_mask_w1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.545 0.070 90.615 ;
    END
  END w_mask_w1[21]
  PIN w_mask_w1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.885 0.070 94.955 ;
    END
  END w_mask_w1[22]
  PIN w_mask_w1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.225 0.070 99.295 ;
    END
  END w_mask_w1[23]
  PIN w_mask_w1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.565 0.070 103.635 ;
    END
  END w_mask_w1[24]
  PIN w_mask_w1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.905 0.070 107.975 ;
    END
  END w_mask_w1[25]
  PIN w_mask_w1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.245 0.070 112.315 ;
    END
  END w_mask_w1[26]
  PIN w_mask_w1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.585 0.070 116.655 ;
    END
  END w_mask_w1[27]
  PIN w_mask_w1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.925 0.070 120.995 ;
    END
  END w_mask_w1[28]
  PIN w_mask_w1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.265 0.070 125.335 ;
    END
  END w_mask_w1[29]
  PIN w_mask_w1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.605 0.070 129.675 ;
    END
  END w_mask_w1[30]
  PIN w_mask_w1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.945 0.070 134.015 ;
    END
  END w_mask_w1[31]
  PIN rd_out_r1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.325 0.070 136.395 ;
    END
  END rd_out_r1[0]
  PIN rd_out_r1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.665 0.070 140.735 ;
    END
  END rd_out_r1[1]
  PIN rd_out_r1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.005 0.070 145.075 ;
    END
  END rd_out_r1[2]
  PIN rd_out_r1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.345 0.070 149.415 ;
    END
  END rd_out_r1[3]
  PIN rd_out_r1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.685 0.070 153.755 ;
    END
  END rd_out_r1[4]
  PIN rd_out_r1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.025 0.070 158.095 ;
    END
  END rd_out_r1[5]
  PIN rd_out_r1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.365 0.070 162.435 ;
    END
  END rd_out_r1[6]
  PIN rd_out_r1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.705 0.070 166.775 ;
    END
  END rd_out_r1[7]
  PIN rd_out_r1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.045 0.070 171.115 ;
    END
  END rd_out_r1[8]
  PIN rd_out_r1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.385 0.070 175.455 ;
    END
  END rd_out_r1[9]
  PIN rd_out_r1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.725 0.070 179.795 ;
    END
  END rd_out_r1[10]
  PIN rd_out_r1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.065 0.070 184.135 ;
    END
  END rd_out_r1[11]
  PIN rd_out_r1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.405 0.070 188.475 ;
    END
  END rd_out_r1[12]
  PIN rd_out_r1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.745 0.070 192.815 ;
    END
  END rd_out_r1[13]
  PIN rd_out_r1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.085 0.070 197.155 ;
    END
  END rd_out_r1[14]
  PIN rd_out_r1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.425 0.070 201.495 ;
    END
  END rd_out_r1[15]
  PIN rd_out_r1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.765 0.070 205.835 ;
    END
  END rd_out_r1[16]
  PIN rd_out_r1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.105 0.070 210.175 ;
    END
  END rd_out_r1[17]
  PIN rd_out_r1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.445 0.070 214.515 ;
    END
  END rd_out_r1[18]
  PIN rd_out_r1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.785 0.070 218.855 ;
    END
  END rd_out_r1[19]
  PIN rd_out_r1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.125 0.070 223.195 ;
    END
  END rd_out_r1[20]
  PIN rd_out_r1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.465 0.070 227.535 ;
    END
  END rd_out_r1[21]
  PIN rd_out_r1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.805 0.070 231.875 ;
    END
  END rd_out_r1[22]
  PIN rd_out_r1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.145 0.070 236.215 ;
    END
  END rd_out_r1[23]
  PIN rd_out_r1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.485 0.070 240.555 ;
    END
  END rd_out_r1[24]
  PIN rd_out_r1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.825 0.070 244.895 ;
    END
  END rd_out_r1[25]
  PIN rd_out_r1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.165 0.070 249.235 ;
    END
  END rd_out_r1[26]
  PIN rd_out_r1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.505 0.070 253.575 ;
    END
  END rd_out_r1[27]
  PIN rd_out_r1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.845 0.070 257.915 ;
    END
  END rd_out_r1[28]
  PIN rd_out_r1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.185 0.070 262.255 ;
    END
  END rd_out_r1[29]
  PIN rd_out_r1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.525 0.070 266.595 ;
    END
  END rd_out_r1[30]
  PIN rd_out_r1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.865 0.070 270.935 ;
    END
  END rd_out_r1[31]
  PIN wd_in_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.245 0.070 273.315 ;
    END
  END wd_in_w1[0]
  PIN wd_in_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.585 0.070 277.655 ;
    END
  END wd_in_w1[1]
  PIN wd_in_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.925 0.070 281.995 ;
    END
  END wd_in_w1[2]
  PIN wd_in_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.265 0.070 286.335 ;
    END
  END wd_in_w1[3]
  PIN wd_in_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.605 0.070 290.675 ;
    END
  END wd_in_w1[4]
  PIN wd_in_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.945 0.070 295.015 ;
    END
  END wd_in_w1[5]
  PIN wd_in_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.285 0.070 299.355 ;
    END
  END wd_in_w1[6]
  PIN wd_in_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.625 0.070 303.695 ;
    END
  END wd_in_w1[7]
  PIN wd_in_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.965 0.070 308.035 ;
    END
  END wd_in_w1[8]
  PIN wd_in_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.305 0.070 312.375 ;
    END
  END wd_in_w1[9]
  PIN wd_in_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.645 0.070 316.715 ;
    END
  END wd_in_w1[10]
  PIN wd_in_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.985 0.070 321.055 ;
    END
  END wd_in_w1[11]
  PIN wd_in_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.325 0.070 325.395 ;
    END
  END wd_in_w1[12]
  PIN wd_in_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.665 0.070 329.735 ;
    END
  END wd_in_w1[13]
  PIN wd_in_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.005 0.070 334.075 ;
    END
  END wd_in_w1[14]
  PIN wd_in_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.345 0.070 338.415 ;
    END
  END wd_in_w1[15]
  PIN wd_in_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.685 0.070 342.755 ;
    END
  END wd_in_w1[16]
  PIN wd_in_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.025 0.070 347.095 ;
    END
  END wd_in_w1[17]
  PIN wd_in_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.365 0.070 351.435 ;
    END
  END wd_in_w1[18]
  PIN wd_in_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.705 0.070 355.775 ;
    END
  END wd_in_w1[19]
  PIN wd_in_w1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.045 0.070 360.115 ;
    END
  END wd_in_w1[20]
  PIN wd_in_w1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.385 0.070 364.455 ;
    END
  END wd_in_w1[21]
  PIN wd_in_w1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.725 0.070 368.795 ;
    END
  END wd_in_w1[22]
  PIN wd_in_w1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.065 0.070 373.135 ;
    END
  END wd_in_w1[23]
  PIN wd_in_w1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.405 0.070 377.475 ;
    END
  END wd_in_w1[24]
  PIN wd_in_w1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.745 0.070 381.815 ;
    END
  END wd_in_w1[25]
  PIN wd_in_w1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.085 0.070 386.155 ;
    END
  END wd_in_w1[26]
  PIN wd_in_w1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.425 0.070 390.495 ;
    END
  END wd_in_w1[27]
  PIN wd_in_w1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.765 0.070 394.835 ;
    END
  END wd_in_w1[28]
  PIN wd_in_w1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.105 0.070 399.175 ;
    END
  END wd_in_w1[29]
  PIN wd_in_w1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 403.445 0.070 403.515 ;
    END
  END wd_in_w1[30]
  PIN wd_in_w1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 407.785 0.070 407.855 ;
    END
  END wd_in_w1[31]
  PIN addr_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 410.165 0.070 410.235 ;
    END
  END addr_w1[0]
  PIN addr_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 414.505 0.070 414.575 ;
    END
  END addr_w1[1]
  PIN addr_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 418.845 0.070 418.915 ;
    END
  END addr_w1[2]
  PIN addr_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 423.185 0.070 423.255 ;
    END
  END addr_w1[3]
  PIN addr_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 427.525 0.070 427.595 ;
    END
  END addr_w1[4]
  PIN addr_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 431.865 0.070 431.935 ;
    END
  END addr_w1[5]
  PIN addr_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 436.205 0.070 436.275 ;
    END
  END addr_w1[6]
  PIN addr_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 440.545 0.070 440.615 ;
    END
  END addr_w1[7]
  PIN addr_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 444.885 0.070 444.955 ;
    END
  END addr_w1[8]
  PIN addr_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 449.225 0.070 449.295 ;
    END
  END addr_w1[9]
  PIN addr_r1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 451.605 0.070 451.675 ;
    END
  END addr_r1[0]
  PIN addr_r1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 455.945 0.070 456.015 ;
    END
  END addr_r1[1]
  PIN addr_r1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 460.285 0.070 460.355 ;
    END
  END addr_r1[2]
  PIN addr_r1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 464.625 0.070 464.695 ;
    END
  END addr_r1[3]
  PIN addr_r1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 468.965 0.070 469.035 ;
    END
  END addr_r1[4]
  PIN addr_r1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 473.305 0.070 473.375 ;
    END
  END addr_r1[5]
  PIN addr_r1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 477.645 0.070 477.715 ;
    END
  END addr_r1[6]
  PIN addr_r1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 481.985 0.070 482.055 ;
    END
  END addr_r1[7]
  PIN addr_r1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 486.325 0.070 486.395 ;
    END
  END addr_r1[8]
  PIN addr_r1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 490.665 0.070 490.735 ;
    END
  END addr_r1[9]
  PIN we_in_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 493.045 0.070 493.115 ;
    END
  END we_in_w1
  PIN ce_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 493.465 0.070 493.535 ;
    END
  END ce_w1
  PIN ce_r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 495.845 0.070 495.915 ;
    END
  END ce_r1
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 498.225 0.070 498.295 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 484.400 ;
      RECT 3.500 1.400 3.780 484.400 ;
      RECT 5.740 1.400 6.020 484.400 ;
      RECT 7.980 1.400 8.260 484.400 ;
      RECT 10.220 1.400 10.500 484.400 ;
      RECT 12.460 1.400 12.740 484.400 ;
      RECT 14.700 1.400 14.980 484.400 ;
      RECT 16.940 1.400 17.220 484.400 ;
      RECT 19.180 1.400 19.460 484.400 ;
      RECT 21.420 1.400 21.700 484.400 ;
      RECT 23.660 1.400 23.940 484.400 ;
      RECT 25.900 1.400 26.180 484.400 ;
      RECT 28.140 1.400 28.420 484.400 ;
      RECT 30.380 1.400 30.660 484.400 ;
      RECT 32.620 1.400 32.900 484.400 ;
      RECT 34.860 1.400 35.140 484.400 ;
      RECT 37.100 1.400 37.380 484.400 ;
      RECT 39.340 1.400 39.620 484.400 ;
      RECT 41.580 1.400 41.860 484.400 ;
      RECT 43.820 1.400 44.100 484.400 ;
      RECT 46.060 1.400 46.340 484.400 ;
      RECT 48.300 1.400 48.580 484.400 ;
      RECT 50.540 1.400 50.820 484.400 ;
      RECT 52.780 1.400 53.060 484.400 ;
      RECT 55.020 1.400 55.300 484.400 ;
      RECT 57.260 1.400 57.540 484.400 ;
      RECT 59.500 1.400 59.780 484.400 ;
      RECT 61.740 1.400 62.020 484.400 ;
      RECT 63.980 1.400 64.260 484.400 ;
      RECT 66.220 1.400 66.500 484.400 ;
      RECT 68.460 1.400 68.740 484.400 ;
      RECT 70.700 1.400 70.980 484.400 ;
      RECT 72.940 1.400 73.220 484.400 ;
      RECT 75.180 1.400 75.460 484.400 ;
      RECT 77.420 1.400 77.700 484.400 ;
      RECT 79.660 1.400 79.940 484.400 ;
      RECT 81.900 1.400 82.180 484.400 ;
      RECT 84.140 1.400 84.420 484.400 ;
      RECT 86.380 1.400 86.660 484.400 ;
      RECT 88.620 1.400 88.900 484.400 ;
      RECT 90.860 1.400 91.140 484.400 ;
      RECT 93.100 1.400 93.380 484.400 ;
      RECT 95.340 1.400 95.620 484.400 ;
      RECT 97.580 1.400 97.860 484.400 ;
      RECT 99.820 1.400 100.100 484.400 ;
      RECT 102.060 1.400 102.340 484.400 ;
      RECT 104.300 1.400 104.580 484.400 ;
      RECT 106.540 1.400 106.820 484.400 ;
      RECT 108.780 1.400 109.060 484.400 ;
      RECT 111.020 1.400 111.300 484.400 ;
      RECT 113.260 1.400 113.540 484.400 ;
      RECT 115.500 1.400 115.780 484.400 ;
      RECT 117.740 1.400 118.020 484.400 ;
      RECT 119.980 1.400 120.260 484.400 ;
      RECT 122.220 1.400 122.500 484.400 ;
      RECT 124.460 1.400 124.740 484.400 ;
      RECT 126.700 1.400 126.980 484.400 ;
      RECT 128.940 1.400 129.220 484.400 ;
      RECT 131.180 1.400 131.460 484.400 ;
      RECT 133.420 1.400 133.700 484.400 ;
      RECT 135.660 1.400 135.940 484.400 ;
      RECT 137.900 1.400 138.180 484.400 ;
      RECT 140.140 1.400 140.420 484.400 ;
      RECT 142.380 1.400 142.660 484.400 ;
      RECT 144.620 1.400 144.900 484.400 ;
      RECT 146.860 1.400 147.140 484.400 ;
      RECT 149.100 1.400 149.380 484.400 ;
      RECT 151.340 1.400 151.620 484.400 ;
      RECT 153.580 1.400 153.860 484.400 ;
      RECT 155.820 1.400 156.100 484.400 ;
      RECT 158.060 1.400 158.340 484.400 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 484.400 ;
      RECT 4.620 1.400 4.900 484.400 ;
      RECT 6.860 1.400 7.140 484.400 ;
      RECT 9.100 1.400 9.380 484.400 ;
      RECT 11.340 1.400 11.620 484.400 ;
      RECT 13.580 1.400 13.860 484.400 ;
      RECT 15.820 1.400 16.100 484.400 ;
      RECT 18.060 1.400 18.340 484.400 ;
      RECT 20.300 1.400 20.580 484.400 ;
      RECT 22.540 1.400 22.820 484.400 ;
      RECT 24.780 1.400 25.060 484.400 ;
      RECT 27.020 1.400 27.300 484.400 ;
      RECT 29.260 1.400 29.540 484.400 ;
      RECT 31.500 1.400 31.780 484.400 ;
      RECT 33.740 1.400 34.020 484.400 ;
      RECT 35.980 1.400 36.260 484.400 ;
      RECT 38.220 1.400 38.500 484.400 ;
      RECT 40.460 1.400 40.740 484.400 ;
      RECT 42.700 1.400 42.980 484.400 ;
      RECT 44.940 1.400 45.220 484.400 ;
      RECT 47.180 1.400 47.460 484.400 ;
      RECT 49.420 1.400 49.700 484.400 ;
      RECT 51.660 1.400 51.940 484.400 ;
      RECT 53.900 1.400 54.180 484.400 ;
      RECT 56.140 1.400 56.420 484.400 ;
      RECT 58.380 1.400 58.660 484.400 ;
      RECT 60.620 1.400 60.900 484.400 ;
      RECT 62.860 1.400 63.140 484.400 ;
      RECT 65.100 1.400 65.380 484.400 ;
      RECT 67.340 1.400 67.620 484.400 ;
      RECT 69.580 1.400 69.860 484.400 ;
      RECT 71.820 1.400 72.100 484.400 ;
      RECT 74.060 1.400 74.340 484.400 ;
      RECT 76.300 1.400 76.580 484.400 ;
      RECT 78.540 1.400 78.820 484.400 ;
      RECT 80.780 1.400 81.060 484.400 ;
      RECT 83.020 1.400 83.300 484.400 ;
      RECT 85.260 1.400 85.540 484.400 ;
      RECT 87.500 1.400 87.780 484.400 ;
      RECT 89.740 1.400 90.020 484.400 ;
      RECT 91.980 1.400 92.260 484.400 ;
      RECT 94.220 1.400 94.500 484.400 ;
      RECT 96.460 1.400 96.740 484.400 ;
      RECT 98.700 1.400 98.980 484.400 ;
      RECT 100.940 1.400 101.220 484.400 ;
      RECT 103.180 1.400 103.460 484.400 ;
      RECT 105.420 1.400 105.700 484.400 ;
      RECT 107.660 1.400 107.940 484.400 ;
      RECT 109.900 1.400 110.180 484.400 ;
      RECT 112.140 1.400 112.420 484.400 ;
      RECT 114.380 1.400 114.660 484.400 ;
      RECT 116.620 1.400 116.900 484.400 ;
      RECT 118.860 1.400 119.140 484.400 ;
      RECT 121.100 1.400 121.380 484.400 ;
      RECT 123.340 1.400 123.620 484.400 ;
      RECT 125.580 1.400 125.860 484.400 ;
      RECT 127.820 1.400 128.100 484.400 ;
      RECT 130.060 1.400 130.340 484.400 ;
      RECT 132.300 1.400 132.580 484.400 ;
      RECT 134.540 1.400 134.820 484.400 ;
      RECT 136.780 1.400 137.060 484.400 ;
      RECT 139.020 1.400 139.300 484.400 ;
      RECT 141.260 1.400 141.540 484.400 ;
      RECT 143.500 1.400 143.780 484.400 ;
      RECT 145.740 1.400 146.020 484.400 ;
      RECT 147.980 1.400 148.260 484.400 ;
      RECT 150.220 1.400 150.500 484.400 ;
      RECT 152.460 1.400 152.740 484.400 ;
      RECT 154.700 1.400 154.980 484.400 ;
      RECT 156.940 1.400 157.220 484.400 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 159.980 485.800 ;
    LAYER metal2 ;
    RECT 0 0 159.980 485.800 ;
    LAYER metal3 ;
    RECT 0.070 0 159.980 485.800 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 5.705 ;
    RECT 0 5.775 0.070 10.045 ;
    RECT 0 10.115 0.070 14.385 ;
    RECT 0 14.455 0.070 18.725 ;
    RECT 0 18.795 0.070 23.065 ;
    RECT 0 23.135 0.070 27.405 ;
    RECT 0 27.475 0.070 31.745 ;
    RECT 0 31.815 0.070 36.085 ;
    RECT 0 36.155 0.070 40.425 ;
    RECT 0 40.495 0.070 44.765 ;
    RECT 0 44.835 0.070 49.105 ;
    RECT 0 49.175 0.070 53.445 ;
    RECT 0 53.515 0.070 57.785 ;
    RECT 0 57.855 0.070 62.125 ;
    RECT 0 62.195 0.070 66.465 ;
    RECT 0 66.535 0.070 70.805 ;
    RECT 0 70.875 0.070 75.145 ;
    RECT 0 75.215 0.070 79.485 ;
    RECT 0 79.555 0.070 83.825 ;
    RECT 0 83.895 0.070 88.165 ;
    RECT 0 88.235 0.070 92.505 ;
    RECT 0 92.575 0.070 96.845 ;
    RECT 0 96.915 0.070 101.185 ;
    RECT 0 101.255 0.070 105.525 ;
    RECT 0 105.595 0.070 109.865 ;
    RECT 0 109.935 0.070 114.205 ;
    RECT 0 114.275 0.070 118.545 ;
    RECT 0 118.615 0.070 122.885 ;
    RECT 0 122.955 0.070 127.225 ;
    RECT 0 127.295 0.070 131.565 ;
    RECT 0 131.635 0.070 135.905 ;
    RECT 0 135.975 0.070 138.285 ;
    RECT 0 138.355 0.070 142.625 ;
    RECT 0 142.695 0.070 146.965 ;
    RECT 0 147.035 0.070 151.305 ;
    RECT 0 151.375 0.070 155.645 ;
    RECT 0 155.715 0.070 159.985 ;
    RECT 0 160.055 0.070 164.325 ;
    RECT 0 164.395 0.070 168.665 ;
    RECT 0 168.735 0.070 173.005 ;
    RECT 0 173.075 0.070 177.345 ;
    RECT 0 177.415 0.070 181.685 ;
    RECT 0 181.755 0.070 186.025 ;
    RECT 0 186.095 0.070 190.365 ;
    RECT 0 190.435 0.070 194.705 ;
    RECT 0 194.775 0.070 199.045 ;
    RECT 0 199.115 0.070 203.385 ;
    RECT 0 203.455 0.070 207.725 ;
    RECT 0 207.795 0.070 212.065 ;
    RECT 0 212.135 0.070 216.405 ;
    RECT 0 216.475 0.070 220.745 ;
    RECT 0 220.815 0.070 225.085 ;
    RECT 0 225.155 0.070 229.425 ;
    RECT 0 229.495 0.070 233.765 ;
    RECT 0 233.835 0.070 238.105 ;
    RECT 0 238.175 0.070 242.445 ;
    RECT 0 242.515 0.070 246.785 ;
    RECT 0 246.855 0.070 251.125 ;
    RECT 0 251.195 0.070 255.465 ;
    RECT 0 255.535 0.070 259.805 ;
    RECT 0 259.875 0.070 264.145 ;
    RECT 0 264.215 0.070 268.485 ;
    RECT 0 268.555 0.070 272.825 ;
    RECT 0 272.895 0.070 275.205 ;
    RECT 0 275.275 0.070 279.545 ;
    RECT 0 279.615 0.070 283.885 ;
    RECT 0 283.955 0.070 288.225 ;
    RECT 0 288.295 0.070 292.565 ;
    RECT 0 292.635 0.070 296.905 ;
    RECT 0 296.975 0.070 301.245 ;
    RECT 0 301.315 0.070 305.585 ;
    RECT 0 305.655 0.070 309.925 ;
    RECT 0 309.995 0.070 314.265 ;
    RECT 0 314.335 0.070 318.605 ;
    RECT 0 318.675 0.070 322.945 ;
    RECT 0 323.015 0.070 327.285 ;
    RECT 0 327.355 0.070 331.625 ;
    RECT 0 331.695 0.070 335.965 ;
    RECT 0 336.035 0.070 340.305 ;
    RECT 0 340.375 0.070 344.645 ;
    RECT 0 344.715 0.070 348.985 ;
    RECT 0 349.055 0.070 353.325 ;
    RECT 0 353.395 0.070 357.665 ;
    RECT 0 357.735 0.070 362.005 ;
    RECT 0 362.075 0.070 366.345 ;
    RECT 0 366.415 0.070 370.685 ;
    RECT 0 370.755 0.070 375.025 ;
    RECT 0 375.095 0.070 379.365 ;
    RECT 0 379.435 0.070 383.705 ;
    RECT 0 383.775 0.070 388.045 ;
    RECT 0 388.115 0.070 392.385 ;
    RECT 0 392.455 0.070 396.725 ;
    RECT 0 396.795 0.070 401.065 ;
    RECT 0 401.135 0.070 405.405 ;
    RECT 0 405.475 0.070 409.745 ;
    RECT 0 409.815 0.070 412.125 ;
    RECT 0 412.195 0.070 416.465 ;
    RECT 0 416.535 0.070 420.805 ;
    RECT 0 420.875 0.070 425.145 ;
    RECT 0 425.215 0.070 429.485 ;
    RECT 0 429.555 0.070 433.825 ;
    RECT 0 433.895 0.070 438.165 ;
    RECT 0 438.235 0.070 442.505 ;
    RECT 0 442.575 0.070 446.845 ;
    RECT 0 446.915 0.070 451.185 ;
    RECT 0 451.255 0.070 453.565 ;
    RECT 0 453.635 0.070 457.905 ;
    RECT 0 457.975 0.070 462.245 ;
    RECT 0 462.315 0.070 485.800 ;
    LAYER metal4 ;
    RECT 0 0 159.980 1.400 ;
    RECT 0 484.400 159.980 485.800 ;
    RECT 0.000 1.400 1.260 484.400 ;
    RECT 1.540 1.400 2.380 484.400 ;
    RECT 2.660 1.400 3.500 484.400 ;
    RECT 3.780 1.400 4.620 484.400 ;
    RECT 4.900 1.400 5.740 484.400 ;
    RECT 6.020 1.400 6.860 484.400 ;
    RECT 7.140 1.400 7.980 484.400 ;
    RECT 8.260 1.400 9.100 484.400 ;
    RECT 9.380 1.400 10.220 484.400 ;
    RECT 10.500 1.400 11.340 484.400 ;
    RECT 11.620 1.400 12.460 484.400 ;
    RECT 12.740 1.400 13.580 484.400 ;
    RECT 13.860 1.400 14.700 484.400 ;
    RECT 14.980 1.400 15.820 484.400 ;
    RECT 16.100 1.400 16.940 484.400 ;
    RECT 17.220 1.400 18.060 484.400 ;
    RECT 18.340 1.400 19.180 484.400 ;
    RECT 19.460 1.400 20.300 484.400 ;
    RECT 20.580 1.400 21.420 484.400 ;
    RECT 21.700 1.400 22.540 484.400 ;
    RECT 22.820 1.400 23.660 484.400 ;
    RECT 23.940 1.400 24.780 484.400 ;
    RECT 25.060 1.400 25.900 484.400 ;
    RECT 26.180 1.400 27.020 484.400 ;
    RECT 27.300 1.400 28.140 484.400 ;
    RECT 28.420 1.400 29.260 484.400 ;
    RECT 29.540 1.400 30.380 484.400 ;
    RECT 30.660 1.400 31.500 484.400 ;
    RECT 31.780 1.400 32.620 484.400 ;
    RECT 32.900 1.400 33.740 484.400 ;
    RECT 34.020 1.400 34.860 484.400 ;
    RECT 35.140 1.400 35.980 484.400 ;
    RECT 36.260 1.400 37.100 484.400 ;
    RECT 37.380 1.400 38.220 484.400 ;
    RECT 38.500 1.400 39.340 484.400 ;
    RECT 39.620 1.400 40.460 484.400 ;
    RECT 40.740 1.400 41.580 484.400 ;
    RECT 41.860 1.400 42.700 484.400 ;
    RECT 42.980 1.400 43.820 484.400 ;
    RECT 44.100 1.400 44.940 484.400 ;
    RECT 45.220 1.400 46.060 484.400 ;
    RECT 46.340 1.400 47.180 484.400 ;
    RECT 47.460 1.400 48.300 484.400 ;
    RECT 48.580 1.400 49.420 484.400 ;
    RECT 49.700 1.400 50.540 484.400 ;
    RECT 50.820 1.400 51.660 484.400 ;
    RECT 51.940 1.400 52.780 484.400 ;
    RECT 53.060 1.400 53.900 484.400 ;
    RECT 54.180 1.400 55.020 484.400 ;
    RECT 55.300 1.400 56.140 484.400 ;
    RECT 56.420 1.400 57.260 484.400 ;
    RECT 57.540 1.400 58.380 484.400 ;
    RECT 58.660 1.400 59.500 484.400 ;
    RECT 59.780 1.400 60.620 484.400 ;
    RECT 60.900 1.400 61.740 484.400 ;
    RECT 62.020 1.400 62.860 484.400 ;
    RECT 63.140 1.400 63.980 484.400 ;
    RECT 64.260 1.400 65.100 484.400 ;
    RECT 65.380 1.400 66.220 484.400 ;
    RECT 66.500 1.400 67.340 484.400 ;
    RECT 67.620 1.400 68.460 484.400 ;
    RECT 68.740 1.400 69.580 484.400 ;
    RECT 69.860 1.400 70.700 484.400 ;
    RECT 70.980 1.400 71.820 484.400 ;
    RECT 72.100 1.400 72.940 484.400 ;
    RECT 73.220 1.400 74.060 484.400 ;
    RECT 74.340 1.400 75.180 484.400 ;
    RECT 75.460 1.400 76.300 484.400 ;
    RECT 76.580 1.400 77.420 484.400 ;
    RECT 77.700 1.400 78.540 484.400 ;
    RECT 78.820 1.400 79.660 484.400 ;
    RECT 79.940 1.400 80.780 484.400 ;
    RECT 81.060 1.400 81.900 484.400 ;
    RECT 82.180 1.400 83.020 484.400 ;
    RECT 83.300 1.400 84.140 484.400 ;
    RECT 84.420 1.400 85.260 484.400 ;
    RECT 85.540 1.400 86.380 484.400 ;
    RECT 86.660 1.400 87.500 484.400 ;
    RECT 87.780 1.400 88.620 484.400 ;
    RECT 88.900 1.400 89.740 484.400 ;
    RECT 90.020 1.400 90.860 484.400 ;
    RECT 91.140 1.400 91.980 484.400 ;
    RECT 92.260 1.400 93.100 484.400 ;
    RECT 93.380 1.400 94.220 484.400 ;
    RECT 94.500 1.400 95.340 484.400 ;
    RECT 95.620 1.400 96.460 484.400 ;
    RECT 96.740 1.400 97.580 484.400 ;
    RECT 97.860 1.400 98.700 484.400 ;
    RECT 98.980 1.400 99.820 484.400 ;
    RECT 100.100 1.400 100.940 484.400 ;
    RECT 101.220 1.400 102.060 484.400 ;
    RECT 102.340 1.400 103.180 484.400 ;
    RECT 103.460 1.400 104.300 484.400 ;
    RECT 104.580 1.400 105.420 484.400 ;
    RECT 105.700 1.400 106.540 484.400 ;
    RECT 106.820 1.400 107.660 484.400 ;
    RECT 107.940 1.400 108.780 484.400 ;
    RECT 109.060 1.400 109.900 484.400 ;
    RECT 110.180 1.400 111.020 484.400 ;
    RECT 111.300 1.400 112.140 484.400 ;
    RECT 112.420 1.400 113.260 484.400 ;
    RECT 113.540 1.400 114.380 484.400 ;
    RECT 114.660 1.400 115.500 484.400 ;
    RECT 115.780 1.400 116.620 484.400 ;
    RECT 116.900 1.400 117.740 484.400 ;
    RECT 118.020 1.400 118.860 484.400 ;
    RECT 119.140 1.400 119.980 484.400 ;
    RECT 120.260 1.400 121.100 484.400 ;
    RECT 121.380 1.400 122.220 484.400 ;
    RECT 122.500 1.400 123.340 484.400 ;
    RECT 123.620 1.400 124.460 484.400 ;
    RECT 124.740 1.400 125.580 484.400 ;
    RECT 125.860 1.400 126.700 484.400 ;
    RECT 126.980 1.400 127.820 484.400 ;
    RECT 128.100 1.400 128.940 484.400 ;
    RECT 129.220 1.400 130.060 484.400 ;
    RECT 130.340 1.400 131.180 484.400 ;
    RECT 131.460 1.400 132.300 484.400 ;
    RECT 132.580 1.400 133.420 484.400 ;
    RECT 133.700 1.400 134.540 484.400 ;
    RECT 134.820 1.400 135.660 484.400 ;
    RECT 135.940 1.400 136.780 484.400 ;
    RECT 137.060 1.400 137.900 484.400 ;
    RECT 138.180 1.400 139.020 484.400 ;
    RECT 139.300 1.400 140.140 484.400 ;
    RECT 140.420 1.400 141.260 484.400 ;
    RECT 141.540 1.400 142.380 484.400 ;
    RECT 142.660 1.400 143.500 484.400 ;
    RECT 143.780 1.400 144.620 484.400 ;
    RECT 144.900 1.400 145.740 484.400 ;
    RECT 146.020 1.400 146.860 484.400 ;
    RECT 147.140 1.400 147.980 484.400 ;
    RECT 148.260 1.400 149.100 484.400 ;
    RECT 149.380 1.400 150.220 484.400 ;
    RECT 150.500 1.400 151.340 484.400 ;
    RECT 151.620 1.400 152.460 484.400 ;
    RECT 152.740 1.400 153.580 484.400 ;
    RECT 153.860 1.400 154.700 484.400 ;
    RECT 154.980 1.400 155.820 484.400 ;
    RECT 156.100 1.400 156.940 484.400 ;
    RECT 157.220 1.400 158.060 484.400 ;
    RECT 158.340 1.400 159.980 484.400 ;
    LAYER OVERLAP ;
    RECT 0 0 159.980 485.800 ;
  END
END sram_32x1024_1r1w

END LIBRARY
