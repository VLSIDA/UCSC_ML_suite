VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_20x64_1r1w
  FOREIGN fakeram_20x64_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 76.950 BY 63.000 ;
  CLASS BLOCK ;
  PIN w_mask_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.085 0.070 1.155 ;
    END
  END w_mask_w1[0]
  PIN w_mask_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.925 0.070 1.995 ;
    END
  END w_mask_w1[1]
  PIN w_mask_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_w1[2]
  PIN w_mask_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.605 0.070 3.675 ;
    END
  END w_mask_w1[3]
  PIN w_mask_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.445 0.070 4.515 ;
    END
  END w_mask_w1[4]
  PIN w_mask_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_w1[5]
  PIN w_mask_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.125 0.070 6.195 ;
    END
  END w_mask_w1[6]
  PIN w_mask_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_w1[7]
  PIN w_mask_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.805 0.070 7.875 ;
    END
  END w_mask_w1[8]
  PIN w_mask_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.645 0.070 8.715 ;
    END
  END w_mask_w1[9]
  PIN w_mask_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.485 0.070 9.555 ;
    END
  END w_mask_w1[10]
  PIN w_mask_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.325 0.070 10.395 ;
    END
  END w_mask_w1[11]
  PIN w_mask_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_w1[12]
  PIN w_mask_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.005 0.070 12.075 ;
    END
  END w_mask_w1[13]
  PIN w_mask_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.845 0.070 12.915 ;
    END
  END w_mask_w1[14]
  PIN w_mask_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.685 0.070 13.755 ;
    END
  END w_mask_w1[15]
  PIN w_mask_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.525 0.070 14.595 ;
    END
  END w_mask_w1[16]
  PIN w_mask_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_w1[17]
  PIN w_mask_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.205 0.070 16.275 ;
    END
  END w_mask_w1[18]
  PIN w_mask_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.045 0.070 17.115 ;
    END
  END w_mask_w1[19]
  PIN rd_out_r1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END rd_out_r1[0]
  PIN rd_out_r1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END rd_out_r1[1]
  PIN rd_out_r1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END rd_out_r1[2]
  PIN rd_out_r1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END rd_out_r1[3]
  PIN rd_out_r1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END rd_out_r1[4]
  PIN rd_out_r1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END rd_out_r1[5]
  PIN rd_out_r1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END rd_out_r1[6]
  PIN rd_out_r1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END rd_out_r1[7]
  PIN rd_out_r1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END rd_out_r1[8]
  PIN rd_out_r1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END rd_out_r1[9]
  PIN rd_out_r1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END rd_out_r1[10]
  PIN rd_out_r1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END rd_out_r1[11]
  PIN rd_out_r1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END rd_out_r1[12]
  PIN rd_out_r1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END rd_out_r1[13]
  PIN rd_out_r1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END rd_out_r1[14]
  PIN rd_out_r1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END rd_out_r1[15]
  PIN rd_out_r1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END rd_out_r1[16]
  PIN rd_out_r1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END rd_out_r1[17]
  PIN rd_out_r1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END rd_out_r1[18]
  PIN rd_out_r1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END rd_out_r1[19]
  PIN wd_in_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.125 0.070 34.195 ;
    END
  END wd_in_w1[0]
  PIN wd_in_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END wd_in_w1[1]
  PIN wd_in_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.805 0.070 35.875 ;
    END
  END wd_in_w1[2]
  PIN wd_in_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END wd_in_w1[3]
  PIN wd_in_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.485 0.070 37.555 ;
    END
  END wd_in_w1[4]
  PIN wd_in_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.325 0.070 38.395 ;
    END
  END wd_in_w1[5]
  PIN wd_in_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END wd_in_w1[6]
  PIN wd_in_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.005 0.070 40.075 ;
    END
  END wd_in_w1[7]
  PIN wd_in_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.845 0.070 40.915 ;
    END
  END wd_in_w1[8]
  PIN wd_in_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.685 0.070 41.755 ;
    END
  END wd_in_w1[9]
  PIN wd_in_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END wd_in_w1[10]
  PIN wd_in_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END wd_in_w1[11]
  PIN wd_in_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.205 0.070 44.275 ;
    END
  END wd_in_w1[12]
  PIN wd_in_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END wd_in_w1[13]
  PIN wd_in_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.885 0.070 45.955 ;
    END
  END wd_in_w1[14]
  PIN wd_in_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.725 0.070 46.795 ;
    END
  END wd_in_w1[15]
  PIN wd_in_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.565 0.070 47.635 ;
    END
  END wd_in_w1[16]
  PIN wd_in_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END wd_in_w1[17]
  PIN wd_in_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.245 0.070 49.315 ;
    END
  END wd_in_w1[18]
  PIN wd_in_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.085 0.070 50.155 ;
    END
  END wd_in_w1[19]
  PIN addr_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.645 0.070 50.715 ;
    END
  END addr_w1[0]
  PIN addr_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.485 0.070 51.555 ;
    END
  END addr_w1[1]
  PIN addr_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.325 0.070 52.395 ;
    END
  END addr_w1[2]
  PIN addr_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.165 0.070 53.235 ;
    END
  END addr_w1[3]
  PIN addr_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.005 0.070 54.075 ;
    END
  END addr_w1[4]
  PIN addr_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.845 0.070 54.915 ;
    END
  END addr_w1[5]
  PIN addr_r1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END addr_r1[0]
  PIN addr_r1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END addr_r1[1]
  PIN addr_r1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END addr_r1[2]
  PIN addr_r1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END addr_r1[3]
  PIN addr_r1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END addr_r1[4]
  PIN addr_r1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END addr_r1[5]
  PIN we_in_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END we_in_w1
  PIN ce_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END ce_w1
  PIN ce_r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.005 0.070 61.075 ;
    END
  END ce_r1
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.565 0.070 61.635 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 61.600 ;
      RECT 3.500 1.400 3.780 61.600 ;
      RECT 5.740 1.400 6.020 61.600 ;
      RECT 7.980 1.400 8.260 61.600 ;
      RECT 10.220 1.400 10.500 61.600 ;
      RECT 12.460 1.400 12.740 61.600 ;
      RECT 14.700 1.400 14.980 61.600 ;
      RECT 16.940 1.400 17.220 61.600 ;
      RECT 19.180 1.400 19.460 61.600 ;
      RECT 21.420 1.400 21.700 61.600 ;
      RECT 23.660 1.400 23.940 61.600 ;
      RECT 25.900 1.400 26.180 61.600 ;
      RECT 28.140 1.400 28.420 61.600 ;
      RECT 30.380 1.400 30.660 61.600 ;
      RECT 32.620 1.400 32.900 61.600 ;
      RECT 34.860 1.400 35.140 61.600 ;
      RECT 37.100 1.400 37.380 61.600 ;
      RECT 39.340 1.400 39.620 61.600 ;
      RECT 41.580 1.400 41.860 61.600 ;
      RECT 43.820 1.400 44.100 61.600 ;
      RECT 46.060 1.400 46.340 61.600 ;
      RECT 48.300 1.400 48.580 61.600 ;
      RECT 50.540 1.400 50.820 61.600 ;
      RECT 52.780 1.400 53.060 61.600 ;
      RECT 55.020 1.400 55.300 61.600 ;
      RECT 57.260 1.400 57.540 61.600 ;
      RECT 59.500 1.400 59.780 61.600 ;
      RECT 61.740 1.400 62.020 61.600 ;
      RECT 63.980 1.400 64.260 61.600 ;
      RECT 66.220 1.400 66.500 61.600 ;
      RECT 68.460 1.400 68.740 61.600 ;
      RECT 70.700 1.400 70.980 61.600 ;
      RECT 72.940 1.400 73.220 61.600 ;
      RECT 75.180 1.400 75.460 61.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 61.600 ;
      RECT 4.620 1.400 4.900 61.600 ;
      RECT 6.860 1.400 7.140 61.600 ;
      RECT 9.100 1.400 9.380 61.600 ;
      RECT 11.340 1.400 11.620 61.600 ;
      RECT 13.580 1.400 13.860 61.600 ;
      RECT 15.820 1.400 16.100 61.600 ;
      RECT 18.060 1.400 18.340 61.600 ;
      RECT 20.300 1.400 20.580 61.600 ;
      RECT 22.540 1.400 22.820 61.600 ;
      RECT 24.780 1.400 25.060 61.600 ;
      RECT 27.020 1.400 27.300 61.600 ;
      RECT 29.260 1.400 29.540 61.600 ;
      RECT 31.500 1.400 31.780 61.600 ;
      RECT 33.740 1.400 34.020 61.600 ;
      RECT 35.980 1.400 36.260 61.600 ;
      RECT 38.220 1.400 38.500 61.600 ;
      RECT 40.460 1.400 40.740 61.600 ;
      RECT 42.700 1.400 42.980 61.600 ;
      RECT 44.940 1.400 45.220 61.600 ;
      RECT 47.180 1.400 47.460 61.600 ;
      RECT 49.420 1.400 49.700 61.600 ;
      RECT 51.660 1.400 51.940 61.600 ;
      RECT 53.900 1.400 54.180 61.600 ;
      RECT 56.140 1.400 56.420 61.600 ;
      RECT 58.380 1.400 58.660 61.600 ;
      RECT 60.620 1.400 60.900 61.600 ;
      RECT 62.860 1.400 63.140 61.600 ;
      RECT 65.100 1.400 65.380 61.600 ;
      RECT 67.340 1.400 67.620 61.600 ;
      RECT 69.580 1.400 69.860 61.600 ;
      RECT 71.820 1.400 72.100 61.600 ;
      RECT 74.060 1.400 74.340 61.600 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 76.950 63.000 ;
    LAYER metal2 ;
    RECT 0 0 76.950 63.000 ;
    LAYER metal3 ;
    RECT 0.070 0 76.950 63.000 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 2.205 ;
    RECT 0 2.275 0.070 3.045 ;
    RECT 0 3.115 0.070 3.885 ;
    RECT 0 3.955 0.070 4.725 ;
    RECT 0 4.795 0.070 5.565 ;
    RECT 0 5.635 0.070 6.405 ;
    RECT 0 6.475 0.070 7.245 ;
    RECT 0 7.315 0.070 8.085 ;
    RECT 0 8.155 0.070 8.925 ;
    RECT 0 8.995 0.070 9.765 ;
    RECT 0 9.835 0.070 10.605 ;
    RECT 0 10.675 0.070 11.445 ;
    RECT 0 11.515 0.070 12.285 ;
    RECT 0 12.355 0.070 13.125 ;
    RECT 0 13.195 0.070 13.965 ;
    RECT 0 14.035 0.070 14.805 ;
    RECT 0 14.875 0.070 15.645 ;
    RECT 0 15.715 0.070 16.485 ;
    RECT 0 16.555 0.070 17.325 ;
    RECT 0 17.395 0.070 17.885 ;
    RECT 0 17.955 0.070 18.725 ;
    RECT 0 18.795 0.070 19.565 ;
    RECT 0 19.635 0.070 20.405 ;
    RECT 0 20.475 0.070 21.245 ;
    RECT 0 21.315 0.070 22.085 ;
    RECT 0 22.155 0.070 22.925 ;
    RECT 0 22.995 0.070 23.765 ;
    RECT 0 23.835 0.070 24.605 ;
    RECT 0 24.675 0.070 25.445 ;
    RECT 0 25.515 0.070 26.285 ;
    RECT 0 26.355 0.070 27.125 ;
    RECT 0 27.195 0.070 27.965 ;
    RECT 0 28.035 0.070 28.805 ;
    RECT 0 28.875 0.070 29.645 ;
    RECT 0 29.715 0.070 30.485 ;
    RECT 0 30.555 0.070 31.325 ;
    RECT 0 31.395 0.070 32.165 ;
    RECT 0 32.235 0.070 33.005 ;
    RECT 0 33.075 0.070 33.845 ;
    RECT 0 33.915 0.070 34.405 ;
    RECT 0 34.475 0.070 35.245 ;
    RECT 0 35.315 0.070 36.085 ;
    RECT 0 36.155 0.070 36.925 ;
    RECT 0 36.995 0.070 37.765 ;
    RECT 0 37.835 0.070 38.605 ;
    RECT 0 38.675 0.070 39.445 ;
    RECT 0 39.515 0.070 40.285 ;
    RECT 0 40.355 0.070 41.125 ;
    RECT 0 41.195 0.070 41.965 ;
    RECT 0 42.035 0.070 42.805 ;
    RECT 0 42.875 0.070 43.645 ;
    RECT 0 43.715 0.070 44.485 ;
    RECT 0 44.555 0.070 45.325 ;
    RECT 0 45.395 0.070 46.165 ;
    RECT 0 46.235 0.070 47.005 ;
    RECT 0 47.075 0.070 47.845 ;
    RECT 0 47.915 0.070 48.685 ;
    RECT 0 48.755 0.070 49.525 ;
    RECT 0 49.595 0.070 50.365 ;
    RECT 0 50.435 0.070 50.925 ;
    RECT 0 50.995 0.070 51.765 ;
    RECT 0 51.835 0.070 52.605 ;
    RECT 0 52.675 0.070 53.445 ;
    RECT 0 53.515 0.070 54.285 ;
    RECT 0 54.355 0.070 55.125 ;
    RECT 0 55.195 0.070 55.685 ;
    RECT 0 55.755 0.070 56.525 ;
    RECT 0 56.595 0.070 57.365 ;
    RECT 0 57.435 0.070 63.000 ;
    LAYER metal4 ;
    RECT 0 0 76.950 1.400 ;
    RECT 0 61.600 76.950 63.000 ;
    RECT 0.000 1.400 1.260 61.600 ;
    RECT 1.540 1.400 2.380 61.600 ;
    RECT 2.660 1.400 3.500 61.600 ;
    RECT 3.780 1.400 4.620 61.600 ;
    RECT 4.900 1.400 5.740 61.600 ;
    RECT 6.020 1.400 6.860 61.600 ;
    RECT 7.140 1.400 7.980 61.600 ;
    RECT 8.260 1.400 9.100 61.600 ;
    RECT 9.380 1.400 10.220 61.600 ;
    RECT 10.500 1.400 11.340 61.600 ;
    RECT 11.620 1.400 12.460 61.600 ;
    RECT 12.740 1.400 13.580 61.600 ;
    RECT 13.860 1.400 14.700 61.600 ;
    RECT 14.980 1.400 15.820 61.600 ;
    RECT 16.100 1.400 16.940 61.600 ;
    RECT 17.220 1.400 18.060 61.600 ;
    RECT 18.340 1.400 19.180 61.600 ;
    RECT 19.460 1.400 20.300 61.600 ;
    RECT 20.580 1.400 21.420 61.600 ;
    RECT 21.700 1.400 22.540 61.600 ;
    RECT 22.820 1.400 23.660 61.600 ;
    RECT 23.940 1.400 24.780 61.600 ;
    RECT 25.060 1.400 25.900 61.600 ;
    RECT 26.180 1.400 27.020 61.600 ;
    RECT 27.300 1.400 28.140 61.600 ;
    RECT 28.420 1.400 29.260 61.600 ;
    RECT 29.540 1.400 30.380 61.600 ;
    RECT 30.660 1.400 31.500 61.600 ;
    RECT 31.780 1.400 32.620 61.600 ;
    RECT 32.900 1.400 33.740 61.600 ;
    RECT 34.020 1.400 34.860 61.600 ;
    RECT 35.140 1.400 35.980 61.600 ;
    RECT 36.260 1.400 37.100 61.600 ;
    RECT 37.380 1.400 38.220 61.600 ;
    RECT 38.500 1.400 39.340 61.600 ;
    RECT 39.620 1.400 40.460 61.600 ;
    RECT 40.740 1.400 41.580 61.600 ;
    RECT 41.860 1.400 42.700 61.600 ;
    RECT 42.980 1.400 43.820 61.600 ;
    RECT 44.100 1.400 44.940 61.600 ;
    RECT 45.220 1.400 46.060 61.600 ;
    RECT 46.340 1.400 47.180 61.600 ;
    RECT 47.460 1.400 48.300 61.600 ;
    RECT 48.580 1.400 49.420 61.600 ;
    RECT 49.700 1.400 50.540 61.600 ;
    RECT 50.820 1.400 51.660 61.600 ;
    RECT 51.940 1.400 52.780 61.600 ;
    RECT 53.060 1.400 53.900 61.600 ;
    RECT 54.180 1.400 55.020 61.600 ;
    RECT 55.300 1.400 56.140 61.600 ;
    RECT 56.420 1.400 57.260 61.600 ;
    RECT 57.540 1.400 58.380 61.600 ;
    RECT 58.660 1.400 59.500 61.600 ;
    RECT 59.780 1.400 60.620 61.600 ;
    RECT 60.900 1.400 61.740 61.600 ;
    RECT 62.020 1.400 62.860 61.600 ;
    RECT 63.140 1.400 63.980 61.600 ;
    RECT 64.260 1.400 65.100 61.600 ;
    RECT 65.380 1.400 66.220 61.600 ;
    RECT 66.500 1.400 67.340 61.600 ;
    RECT 67.620 1.400 68.460 61.600 ;
    RECT 68.740 1.400 69.580 61.600 ;
    RECT 69.860 1.400 70.700 61.600 ;
    RECT 70.980 1.400 71.820 61.600 ;
    RECT 72.100 1.400 72.940 61.600 ;
    RECT 73.220 1.400 74.060 61.600 ;
    RECT 74.340 1.400 75.180 61.600 ;
    RECT 75.460 1.400 76.950 61.600 ;
    LAYER OVERLAP ;
    RECT 0 0 76.950 63.000 ;
  END
END fakeram_20x64_1r1w

END LIBRARY
