VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_512x1024_1r1w
  FOREIGN sram_512x1024_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 1832.740 BY 981.400 ;
  CLASS BLOCK ;
  PIN w_mask_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END w_mask_w1[0]
  PIN w_mask_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.085 0.070 29.155 ;
    END
  END w_mask_w1[1]
  PIN w_mask_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.645 0.070 29.715 ;
    END
  END w_mask_w1[2]
  PIN w_mask_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END w_mask_w1[3]
  PIN w_mask_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_w1[4]
  PIN w_mask_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.325 0.070 31.395 ;
    END
  END w_mask_w1[5]
  PIN w_mask_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END w_mask_w1[6]
  PIN w_mask_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.445 0.070 32.515 ;
    END
  END w_mask_w1[7]
  PIN w_mask_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.005 0.070 33.075 ;
    END
  END w_mask_w1[8]
  PIN w_mask_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END w_mask_w1[9]
  PIN w_mask_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.125 0.070 34.195 ;
    END
  END w_mask_w1[10]
  PIN w_mask_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.685 0.070 34.755 ;
    END
  END w_mask_w1[11]
  PIN w_mask_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END w_mask_w1[12]
  PIN w_mask_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.805 0.070 35.875 ;
    END
  END w_mask_w1[13]
  PIN w_mask_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.365 0.070 36.435 ;
    END
  END w_mask_w1[14]
  PIN w_mask_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END w_mask_w1[15]
  PIN w_mask_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.485 0.070 37.555 ;
    END
  END w_mask_w1[16]
  PIN w_mask_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.045 0.070 38.115 ;
    END
  END w_mask_w1[17]
  PIN w_mask_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END w_mask_w1[18]
  PIN w_mask_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END w_mask_w1[19]
  PIN w_mask_w1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.725 0.070 39.795 ;
    END
  END w_mask_w1[20]
  PIN w_mask_w1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END w_mask_w1[21]
  PIN w_mask_w1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.845 0.070 40.915 ;
    END
  END w_mask_w1[22]
  PIN w_mask_w1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.405 0.070 41.475 ;
    END
  END w_mask_w1[23]
  PIN w_mask_w1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END w_mask_w1[24]
  PIN w_mask_w1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END w_mask_w1[25]
  PIN w_mask_w1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.085 0.070 43.155 ;
    END
  END w_mask_w1[26]
  PIN w_mask_w1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END w_mask_w1[27]
  PIN w_mask_w1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.205 0.070 44.275 ;
    END
  END w_mask_w1[28]
  PIN w_mask_w1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.765 0.070 44.835 ;
    END
  END w_mask_w1[29]
  PIN w_mask_w1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END w_mask_w1[30]
  PIN w_mask_w1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.885 0.070 45.955 ;
    END
  END w_mask_w1[31]
  PIN w_mask_w1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.445 0.070 46.515 ;
    END
  END w_mask_w1[32]
  PIN w_mask_w1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END w_mask_w1[33]
  PIN w_mask_w1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.565 0.070 47.635 ;
    END
  END w_mask_w1[34]
  PIN w_mask_w1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.125 0.070 48.195 ;
    END
  END w_mask_w1[35]
  PIN w_mask_w1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END w_mask_w1[36]
  PIN w_mask_w1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.245 0.070 49.315 ;
    END
  END w_mask_w1[37]
  PIN w_mask_w1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.805 0.070 49.875 ;
    END
  END w_mask_w1[38]
  PIN w_mask_w1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END w_mask_w1[39]
  PIN w_mask_w1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.925 0.070 50.995 ;
    END
  END w_mask_w1[40]
  PIN w_mask_w1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.485 0.070 51.555 ;
    END
  END w_mask_w1[41]
  PIN w_mask_w1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END w_mask_w1[42]
  PIN w_mask_w1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.605 0.070 52.675 ;
    END
  END w_mask_w1[43]
  PIN w_mask_w1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.165 0.070 53.235 ;
    END
  END w_mask_w1[44]
  PIN w_mask_w1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END w_mask_w1[45]
  PIN w_mask_w1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.285 0.070 54.355 ;
    END
  END w_mask_w1[46]
  PIN w_mask_w1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.845 0.070 54.915 ;
    END
  END w_mask_w1[47]
  PIN w_mask_w1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END w_mask_w1[48]
  PIN w_mask_w1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.965 0.070 56.035 ;
    END
  END w_mask_w1[49]
  PIN w_mask_w1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.525 0.070 56.595 ;
    END
  END w_mask_w1[50]
  PIN w_mask_w1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END w_mask_w1[51]
  PIN w_mask_w1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.645 0.070 57.715 ;
    END
  END w_mask_w1[52]
  PIN w_mask_w1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.205 0.070 58.275 ;
    END
  END w_mask_w1[53]
  PIN w_mask_w1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END w_mask_w1[54]
  PIN w_mask_w1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.325 0.070 59.395 ;
    END
  END w_mask_w1[55]
  PIN w_mask_w1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.885 0.070 59.955 ;
    END
  END w_mask_w1[56]
  PIN w_mask_w1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END w_mask_w1[57]
  PIN w_mask_w1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.005 0.070 61.075 ;
    END
  END w_mask_w1[58]
  PIN w_mask_w1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.565 0.070 61.635 ;
    END
  END w_mask_w1[59]
  PIN w_mask_w1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END w_mask_w1[60]
  PIN w_mask_w1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.685 0.070 62.755 ;
    END
  END w_mask_w1[61]
  PIN w_mask_w1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.245 0.070 63.315 ;
    END
  END w_mask_w1[62]
  PIN w_mask_w1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.805 0.070 63.875 ;
    END
  END w_mask_w1[63]
  PIN w_mask_w1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.365 0.070 64.435 ;
    END
  END w_mask_w1[64]
  PIN w_mask_w1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.925 0.070 64.995 ;
    END
  END w_mask_w1[65]
  PIN w_mask_w1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.485 0.070 65.555 ;
    END
  END w_mask_w1[66]
  PIN w_mask_w1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.045 0.070 66.115 ;
    END
  END w_mask_w1[67]
  PIN w_mask_w1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.605 0.070 66.675 ;
    END
  END w_mask_w1[68]
  PIN w_mask_w1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END w_mask_w1[69]
  PIN w_mask_w1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.725 0.070 67.795 ;
    END
  END w_mask_w1[70]
  PIN w_mask_w1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.285 0.070 68.355 ;
    END
  END w_mask_w1[71]
  PIN w_mask_w1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END w_mask_w1[72]
  PIN w_mask_w1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.405 0.070 69.475 ;
    END
  END w_mask_w1[73]
  PIN w_mask_w1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.965 0.070 70.035 ;
    END
  END w_mask_w1[74]
  PIN w_mask_w1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END w_mask_w1[75]
  PIN w_mask_w1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.085 0.070 71.155 ;
    END
  END w_mask_w1[76]
  PIN w_mask_w1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.645 0.070 71.715 ;
    END
  END w_mask_w1[77]
  PIN w_mask_w1[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END w_mask_w1[78]
  PIN w_mask_w1[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.765 0.070 72.835 ;
    END
  END w_mask_w1[79]
  PIN w_mask_w1[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.325 0.070 73.395 ;
    END
  END w_mask_w1[80]
  PIN w_mask_w1[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END w_mask_w1[81]
  PIN w_mask_w1[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.445 0.070 74.515 ;
    END
  END w_mask_w1[82]
  PIN w_mask_w1[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.005 0.070 75.075 ;
    END
  END w_mask_w1[83]
  PIN w_mask_w1[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END w_mask_w1[84]
  PIN w_mask_w1[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.125 0.070 76.195 ;
    END
  END w_mask_w1[85]
  PIN w_mask_w1[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.685 0.070 76.755 ;
    END
  END w_mask_w1[86]
  PIN w_mask_w1[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END w_mask_w1[87]
  PIN w_mask_w1[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END w_mask_w1[88]
  PIN w_mask_w1[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.365 0.070 78.435 ;
    END
  END w_mask_w1[89]
  PIN w_mask_w1[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END w_mask_w1[90]
  PIN w_mask_w1[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.485 0.070 79.555 ;
    END
  END w_mask_w1[91]
  PIN w_mask_w1[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.045 0.070 80.115 ;
    END
  END w_mask_w1[92]
  PIN w_mask_w1[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END w_mask_w1[93]
  PIN w_mask_w1[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.165 0.070 81.235 ;
    END
  END w_mask_w1[94]
  PIN w_mask_w1[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.725 0.070 81.795 ;
    END
  END w_mask_w1[95]
  PIN w_mask_w1[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END w_mask_w1[96]
  PIN w_mask_w1[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.845 0.070 82.915 ;
    END
  END w_mask_w1[97]
  PIN w_mask_w1[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.405 0.070 83.475 ;
    END
  END w_mask_w1[98]
  PIN w_mask_w1[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END w_mask_w1[99]
  PIN w_mask_w1[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.525 0.070 84.595 ;
    END
  END w_mask_w1[100]
  PIN w_mask_w1[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.085 0.070 85.155 ;
    END
  END w_mask_w1[101]
  PIN w_mask_w1[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END w_mask_w1[102]
  PIN w_mask_w1[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.205 0.070 86.275 ;
    END
  END w_mask_w1[103]
  PIN w_mask_w1[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.765 0.070 86.835 ;
    END
  END w_mask_w1[104]
  PIN w_mask_w1[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END w_mask_w1[105]
  PIN w_mask_w1[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.885 0.070 87.955 ;
    END
  END w_mask_w1[106]
  PIN w_mask_w1[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.445 0.070 88.515 ;
    END
  END w_mask_w1[107]
  PIN w_mask_w1[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.005 0.070 89.075 ;
    END
  END w_mask_w1[108]
  PIN w_mask_w1[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.565 0.070 89.635 ;
    END
  END w_mask_w1[109]
  PIN w_mask_w1[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.125 0.070 90.195 ;
    END
  END w_mask_w1[110]
  PIN w_mask_w1[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END w_mask_w1[111]
  PIN w_mask_w1[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.245 0.070 91.315 ;
    END
  END w_mask_w1[112]
  PIN w_mask_w1[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.805 0.070 91.875 ;
    END
  END w_mask_w1[113]
  PIN w_mask_w1[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END w_mask_w1[114]
  PIN w_mask_w1[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.925 0.070 92.995 ;
    END
  END w_mask_w1[115]
  PIN w_mask_w1[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.485 0.070 93.555 ;
    END
  END w_mask_w1[116]
  PIN w_mask_w1[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.045 0.070 94.115 ;
    END
  END w_mask_w1[117]
  PIN w_mask_w1[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.605 0.070 94.675 ;
    END
  END w_mask_w1[118]
  PIN w_mask_w1[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.165 0.070 95.235 ;
    END
  END w_mask_w1[119]
  PIN w_mask_w1[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.725 0.070 95.795 ;
    END
  END w_mask_w1[120]
  PIN w_mask_w1[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.285 0.070 96.355 ;
    END
  END w_mask_w1[121]
  PIN w_mask_w1[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.845 0.070 96.915 ;
    END
  END w_mask_w1[122]
  PIN w_mask_w1[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END w_mask_w1[123]
  PIN w_mask_w1[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.965 0.070 98.035 ;
    END
  END w_mask_w1[124]
  PIN w_mask_w1[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.525 0.070 98.595 ;
    END
  END w_mask_w1[125]
  PIN w_mask_w1[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.085 0.070 99.155 ;
    END
  END w_mask_w1[126]
  PIN w_mask_w1[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.645 0.070 99.715 ;
    END
  END w_mask_w1[127]
  PIN w_mask_w1[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.205 0.070 100.275 ;
    END
  END w_mask_w1[128]
  PIN w_mask_w1[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.765 0.070 100.835 ;
    END
  END w_mask_w1[129]
  PIN w_mask_w1[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.325 0.070 101.395 ;
    END
  END w_mask_w1[130]
  PIN w_mask_w1[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.885 0.070 101.955 ;
    END
  END w_mask_w1[131]
  PIN w_mask_w1[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.445 0.070 102.515 ;
    END
  END w_mask_w1[132]
  PIN w_mask_w1[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.005 0.070 103.075 ;
    END
  END w_mask_w1[133]
  PIN w_mask_w1[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.565 0.070 103.635 ;
    END
  END w_mask_w1[134]
  PIN w_mask_w1[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.125 0.070 104.195 ;
    END
  END w_mask_w1[135]
  PIN w_mask_w1[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.685 0.070 104.755 ;
    END
  END w_mask_w1[136]
  PIN w_mask_w1[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.245 0.070 105.315 ;
    END
  END w_mask_w1[137]
  PIN w_mask_w1[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.805 0.070 105.875 ;
    END
  END w_mask_w1[138]
  PIN w_mask_w1[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.365 0.070 106.435 ;
    END
  END w_mask_w1[139]
  PIN w_mask_w1[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.925 0.070 106.995 ;
    END
  END w_mask_w1[140]
  PIN w_mask_w1[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.485 0.070 107.555 ;
    END
  END w_mask_w1[141]
  PIN w_mask_w1[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.045 0.070 108.115 ;
    END
  END w_mask_w1[142]
  PIN w_mask_w1[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.605 0.070 108.675 ;
    END
  END w_mask_w1[143]
  PIN w_mask_w1[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END w_mask_w1[144]
  PIN w_mask_w1[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.725 0.070 109.795 ;
    END
  END w_mask_w1[145]
  PIN w_mask_w1[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.285 0.070 110.355 ;
    END
  END w_mask_w1[146]
  PIN w_mask_w1[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.845 0.070 110.915 ;
    END
  END w_mask_w1[147]
  PIN w_mask_w1[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.405 0.070 111.475 ;
    END
  END w_mask_w1[148]
  PIN w_mask_w1[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.965 0.070 112.035 ;
    END
  END w_mask_w1[149]
  PIN w_mask_w1[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.525 0.070 112.595 ;
    END
  END w_mask_w1[150]
  PIN w_mask_w1[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.085 0.070 113.155 ;
    END
  END w_mask_w1[151]
  PIN w_mask_w1[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.645 0.070 113.715 ;
    END
  END w_mask_w1[152]
  PIN w_mask_w1[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.205 0.070 114.275 ;
    END
  END w_mask_w1[153]
  PIN w_mask_w1[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.765 0.070 114.835 ;
    END
  END w_mask_w1[154]
  PIN w_mask_w1[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.325 0.070 115.395 ;
    END
  END w_mask_w1[155]
  PIN w_mask_w1[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.885 0.070 115.955 ;
    END
  END w_mask_w1[156]
  PIN w_mask_w1[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.445 0.070 116.515 ;
    END
  END w_mask_w1[157]
  PIN w_mask_w1[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.005 0.070 117.075 ;
    END
  END w_mask_w1[158]
  PIN w_mask_w1[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.565 0.070 117.635 ;
    END
  END w_mask_w1[159]
  PIN w_mask_w1[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.125 0.070 118.195 ;
    END
  END w_mask_w1[160]
  PIN w_mask_w1[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.685 0.070 118.755 ;
    END
  END w_mask_w1[161]
  PIN w_mask_w1[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.245 0.070 119.315 ;
    END
  END w_mask_w1[162]
  PIN w_mask_w1[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.805 0.070 119.875 ;
    END
  END w_mask_w1[163]
  PIN w_mask_w1[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.365 0.070 120.435 ;
    END
  END w_mask_w1[164]
  PIN w_mask_w1[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.925 0.070 120.995 ;
    END
  END w_mask_w1[165]
  PIN w_mask_w1[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.485 0.070 121.555 ;
    END
  END w_mask_w1[166]
  PIN w_mask_w1[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.045 0.070 122.115 ;
    END
  END w_mask_w1[167]
  PIN w_mask_w1[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.605 0.070 122.675 ;
    END
  END w_mask_w1[168]
  PIN w_mask_w1[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.165 0.070 123.235 ;
    END
  END w_mask_w1[169]
  PIN w_mask_w1[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.725 0.070 123.795 ;
    END
  END w_mask_w1[170]
  PIN w_mask_w1[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.285 0.070 124.355 ;
    END
  END w_mask_w1[171]
  PIN w_mask_w1[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.845 0.070 124.915 ;
    END
  END w_mask_w1[172]
  PIN w_mask_w1[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.405 0.070 125.475 ;
    END
  END w_mask_w1[173]
  PIN w_mask_w1[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.965 0.070 126.035 ;
    END
  END w_mask_w1[174]
  PIN w_mask_w1[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.525 0.070 126.595 ;
    END
  END w_mask_w1[175]
  PIN w_mask_w1[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.085 0.070 127.155 ;
    END
  END w_mask_w1[176]
  PIN w_mask_w1[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.645 0.070 127.715 ;
    END
  END w_mask_w1[177]
  PIN w_mask_w1[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.205 0.070 128.275 ;
    END
  END w_mask_w1[178]
  PIN w_mask_w1[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.765 0.070 128.835 ;
    END
  END w_mask_w1[179]
  PIN w_mask_w1[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.325 0.070 129.395 ;
    END
  END w_mask_w1[180]
  PIN w_mask_w1[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.885 0.070 129.955 ;
    END
  END w_mask_w1[181]
  PIN w_mask_w1[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.445 0.070 130.515 ;
    END
  END w_mask_w1[182]
  PIN w_mask_w1[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.005 0.070 131.075 ;
    END
  END w_mask_w1[183]
  PIN w_mask_w1[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.565 0.070 131.635 ;
    END
  END w_mask_w1[184]
  PIN w_mask_w1[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.125 0.070 132.195 ;
    END
  END w_mask_w1[185]
  PIN w_mask_w1[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.685 0.070 132.755 ;
    END
  END w_mask_w1[186]
  PIN w_mask_w1[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.245 0.070 133.315 ;
    END
  END w_mask_w1[187]
  PIN w_mask_w1[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.805 0.070 133.875 ;
    END
  END w_mask_w1[188]
  PIN w_mask_w1[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.365 0.070 134.435 ;
    END
  END w_mask_w1[189]
  PIN w_mask_w1[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.925 0.070 134.995 ;
    END
  END w_mask_w1[190]
  PIN w_mask_w1[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.485 0.070 135.555 ;
    END
  END w_mask_w1[191]
  PIN w_mask_w1[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.045 0.070 136.115 ;
    END
  END w_mask_w1[192]
  PIN w_mask_w1[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.605 0.070 136.675 ;
    END
  END w_mask_w1[193]
  PIN w_mask_w1[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.165 0.070 137.235 ;
    END
  END w_mask_w1[194]
  PIN w_mask_w1[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.725 0.070 137.795 ;
    END
  END w_mask_w1[195]
  PIN w_mask_w1[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.285 0.070 138.355 ;
    END
  END w_mask_w1[196]
  PIN w_mask_w1[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.845 0.070 138.915 ;
    END
  END w_mask_w1[197]
  PIN w_mask_w1[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.405 0.070 139.475 ;
    END
  END w_mask_w1[198]
  PIN w_mask_w1[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.965 0.070 140.035 ;
    END
  END w_mask_w1[199]
  PIN w_mask_w1[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.525 0.070 140.595 ;
    END
  END w_mask_w1[200]
  PIN w_mask_w1[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.085 0.070 141.155 ;
    END
  END w_mask_w1[201]
  PIN w_mask_w1[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.645 0.070 141.715 ;
    END
  END w_mask_w1[202]
  PIN w_mask_w1[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.205 0.070 142.275 ;
    END
  END w_mask_w1[203]
  PIN w_mask_w1[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.765 0.070 142.835 ;
    END
  END w_mask_w1[204]
  PIN w_mask_w1[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.325 0.070 143.395 ;
    END
  END w_mask_w1[205]
  PIN w_mask_w1[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.885 0.070 143.955 ;
    END
  END w_mask_w1[206]
  PIN w_mask_w1[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.445 0.070 144.515 ;
    END
  END w_mask_w1[207]
  PIN w_mask_w1[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.005 0.070 145.075 ;
    END
  END w_mask_w1[208]
  PIN w_mask_w1[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.565 0.070 145.635 ;
    END
  END w_mask_w1[209]
  PIN w_mask_w1[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.125 0.070 146.195 ;
    END
  END w_mask_w1[210]
  PIN w_mask_w1[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.685 0.070 146.755 ;
    END
  END w_mask_w1[211]
  PIN w_mask_w1[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.245 0.070 147.315 ;
    END
  END w_mask_w1[212]
  PIN w_mask_w1[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.805 0.070 147.875 ;
    END
  END w_mask_w1[213]
  PIN w_mask_w1[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.365 0.070 148.435 ;
    END
  END w_mask_w1[214]
  PIN w_mask_w1[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.925 0.070 148.995 ;
    END
  END w_mask_w1[215]
  PIN w_mask_w1[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.485 0.070 149.555 ;
    END
  END w_mask_w1[216]
  PIN w_mask_w1[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.045 0.070 150.115 ;
    END
  END w_mask_w1[217]
  PIN w_mask_w1[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.605 0.070 150.675 ;
    END
  END w_mask_w1[218]
  PIN w_mask_w1[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.165 0.070 151.235 ;
    END
  END w_mask_w1[219]
  PIN w_mask_w1[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.725 0.070 151.795 ;
    END
  END w_mask_w1[220]
  PIN w_mask_w1[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.285 0.070 152.355 ;
    END
  END w_mask_w1[221]
  PIN w_mask_w1[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.845 0.070 152.915 ;
    END
  END w_mask_w1[222]
  PIN w_mask_w1[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.405 0.070 153.475 ;
    END
  END w_mask_w1[223]
  PIN w_mask_w1[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.965 0.070 154.035 ;
    END
  END w_mask_w1[224]
  PIN w_mask_w1[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.525 0.070 154.595 ;
    END
  END w_mask_w1[225]
  PIN w_mask_w1[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.085 0.070 155.155 ;
    END
  END w_mask_w1[226]
  PIN w_mask_w1[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.645 0.070 155.715 ;
    END
  END w_mask_w1[227]
  PIN w_mask_w1[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.205 0.070 156.275 ;
    END
  END w_mask_w1[228]
  PIN w_mask_w1[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.765 0.070 156.835 ;
    END
  END w_mask_w1[229]
  PIN w_mask_w1[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.325 0.070 157.395 ;
    END
  END w_mask_w1[230]
  PIN w_mask_w1[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.885 0.070 157.955 ;
    END
  END w_mask_w1[231]
  PIN w_mask_w1[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.445 0.070 158.515 ;
    END
  END w_mask_w1[232]
  PIN w_mask_w1[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.005 0.070 159.075 ;
    END
  END w_mask_w1[233]
  PIN w_mask_w1[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.565 0.070 159.635 ;
    END
  END w_mask_w1[234]
  PIN w_mask_w1[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.125 0.070 160.195 ;
    END
  END w_mask_w1[235]
  PIN w_mask_w1[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.685 0.070 160.755 ;
    END
  END w_mask_w1[236]
  PIN w_mask_w1[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.245 0.070 161.315 ;
    END
  END w_mask_w1[237]
  PIN w_mask_w1[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.805 0.070 161.875 ;
    END
  END w_mask_w1[238]
  PIN w_mask_w1[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.365 0.070 162.435 ;
    END
  END w_mask_w1[239]
  PIN w_mask_w1[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.925 0.070 162.995 ;
    END
  END w_mask_w1[240]
  PIN w_mask_w1[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.485 0.070 163.555 ;
    END
  END w_mask_w1[241]
  PIN w_mask_w1[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.045 0.070 164.115 ;
    END
  END w_mask_w1[242]
  PIN w_mask_w1[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.605 0.070 164.675 ;
    END
  END w_mask_w1[243]
  PIN w_mask_w1[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.165 0.070 165.235 ;
    END
  END w_mask_w1[244]
  PIN w_mask_w1[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.725 0.070 165.795 ;
    END
  END w_mask_w1[245]
  PIN w_mask_w1[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.285 0.070 166.355 ;
    END
  END w_mask_w1[246]
  PIN w_mask_w1[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.845 0.070 166.915 ;
    END
  END w_mask_w1[247]
  PIN w_mask_w1[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.405 0.070 167.475 ;
    END
  END w_mask_w1[248]
  PIN w_mask_w1[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.965 0.070 168.035 ;
    END
  END w_mask_w1[249]
  PIN w_mask_w1[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.525 0.070 168.595 ;
    END
  END w_mask_w1[250]
  PIN w_mask_w1[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.085 0.070 169.155 ;
    END
  END w_mask_w1[251]
  PIN w_mask_w1[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.645 0.070 169.715 ;
    END
  END w_mask_w1[252]
  PIN w_mask_w1[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.205 0.070 170.275 ;
    END
  END w_mask_w1[253]
  PIN w_mask_w1[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.765 0.070 170.835 ;
    END
  END w_mask_w1[254]
  PIN w_mask_w1[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.325 0.070 171.395 ;
    END
  END w_mask_w1[255]
  PIN w_mask_w1[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.885 0.070 171.955 ;
    END
  END w_mask_w1[256]
  PIN w_mask_w1[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.445 0.070 172.515 ;
    END
  END w_mask_w1[257]
  PIN w_mask_w1[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.005 0.070 173.075 ;
    END
  END w_mask_w1[258]
  PIN w_mask_w1[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.565 0.070 173.635 ;
    END
  END w_mask_w1[259]
  PIN w_mask_w1[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.125 0.070 174.195 ;
    END
  END w_mask_w1[260]
  PIN w_mask_w1[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.685 0.070 174.755 ;
    END
  END w_mask_w1[261]
  PIN w_mask_w1[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.245 0.070 175.315 ;
    END
  END w_mask_w1[262]
  PIN w_mask_w1[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.805 0.070 175.875 ;
    END
  END w_mask_w1[263]
  PIN w_mask_w1[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.365 0.070 176.435 ;
    END
  END w_mask_w1[264]
  PIN w_mask_w1[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.925 0.070 176.995 ;
    END
  END w_mask_w1[265]
  PIN w_mask_w1[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.485 0.070 177.555 ;
    END
  END w_mask_w1[266]
  PIN w_mask_w1[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.045 0.070 178.115 ;
    END
  END w_mask_w1[267]
  PIN w_mask_w1[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.605 0.070 178.675 ;
    END
  END w_mask_w1[268]
  PIN w_mask_w1[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.165 0.070 179.235 ;
    END
  END w_mask_w1[269]
  PIN w_mask_w1[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.725 0.070 179.795 ;
    END
  END w_mask_w1[270]
  PIN w_mask_w1[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.285 0.070 180.355 ;
    END
  END w_mask_w1[271]
  PIN w_mask_w1[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.845 0.070 180.915 ;
    END
  END w_mask_w1[272]
  PIN w_mask_w1[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.405 0.070 181.475 ;
    END
  END w_mask_w1[273]
  PIN w_mask_w1[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.965 0.070 182.035 ;
    END
  END w_mask_w1[274]
  PIN w_mask_w1[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.525 0.070 182.595 ;
    END
  END w_mask_w1[275]
  PIN w_mask_w1[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.085 0.070 183.155 ;
    END
  END w_mask_w1[276]
  PIN w_mask_w1[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.645 0.070 183.715 ;
    END
  END w_mask_w1[277]
  PIN w_mask_w1[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.205 0.070 184.275 ;
    END
  END w_mask_w1[278]
  PIN w_mask_w1[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.765 0.070 184.835 ;
    END
  END w_mask_w1[279]
  PIN w_mask_w1[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.325 0.070 185.395 ;
    END
  END w_mask_w1[280]
  PIN w_mask_w1[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.885 0.070 185.955 ;
    END
  END w_mask_w1[281]
  PIN w_mask_w1[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.445 0.070 186.515 ;
    END
  END w_mask_w1[282]
  PIN w_mask_w1[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.005 0.070 187.075 ;
    END
  END w_mask_w1[283]
  PIN w_mask_w1[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.565 0.070 187.635 ;
    END
  END w_mask_w1[284]
  PIN w_mask_w1[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.125 0.070 188.195 ;
    END
  END w_mask_w1[285]
  PIN w_mask_w1[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.685 0.070 188.755 ;
    END
  END w_mask_w1[286]
  PIN w_mask_w1[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.245 0.070 189.315 ;
    END
  END w_mask_w1[287]
  PIN w_mask_w1[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.805 0.070 189.875 ;
    END
  END w_mask_w1[288]
  PIN w_mask_w1[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.365 0.070 190.435 ;
    END
  END w_mask_w1[289]
  PIN w_mask_w1[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.925 0.070 190.995 ;
    END
  END w_mask_w1[290]
  PIN w_mask_w1[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.485 0.070 191.555 ;
    END
  END w_mask_w1[291]
  PIN w_mask_w1[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.045 0.070 192.115 ;
    END
  END w_mask_w1[292]
  PIN w_mask_w1[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.605 0.070 192.675 ;
    END
  END w_mask_w1[293]
  PIN w_mask_w1[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.165 0.070 193.235 ;
    END
  END w_mask_w1[294]
  PIN w_mask_w1[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.725 0.070 193.795 ;
    END
  END w_mask_w1[295]
  PIN w_mask_w1[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.285 0.070 194.355 ;
    END
  END w_mask_w1[296]
  PIN w_mask_w1[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.845 0.070 194.915 ;
    END
  END w_mask_w1[297]
  PIN w_mask_w1[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.405 0.070 195.475 ;
    END
  END w_mask_w1[298]
  PIN w_mask_w1[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.965 0.070 196.035 ;
    END
  END w_mask_w1[299]
  PIN w_mask_w1[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.525 0.070 196.595 ;
    END
  END w_mask_w1[300]
  PIN w_mask_w1[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.085 0.070 197.155 ;
    END
  END w_mask_w1[301]
  PIN w_mask_w1[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.645 0.070 197.715 ;
    END
  END w_mask_w1[302]
  PIN w_mask_w1[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.205 0.070 198.275 ;
    END
  END w_mask_w1[303]
  PIN w_mask_w1[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.765 0.070 198.835 ;
    END
  END w_mask_w1[304]
  PIN w_mask_w1[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.325 0.070 199.395 ;
    END
  END w_mask_w1[305]
  PIN w_mask_w1[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.885 0.070 199.955 ;
    END
  END w_mask_w1[306]
  PIN w_mask_w1[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.445 0.070 200.515 ;
    END
  END w_mask_w1[307]
  PIN w_mask_w1[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.005 0.070 201.075 ;
    END
  END w_mask_w1[308]
  PIN w_mask_w1[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.565 0.070 201.635 ;
    END
  END w_mask_w1[309]
  PIN w_mask_w1[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.125 0.070 202.195 ;
    END
  END w_mask_w1[310]
  PIN w_mask_w1[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.685 0.070 202.755 ;
    END
  END w_mask_w1[311]
  PIN w_mask_w1[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.245 0.070 203.315 ;
    END
  END w_mask_w1[312]
  PIN w_mask_w1[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.805 0.070 203.875 ;
    END
  END w_mask_w1[313]
  PIN w_mask_w1[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.365 0.070 204.435 ;
    END
  END w_mask_w1[314]
  PIN w_mask_w1[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.925 0.070 204.995 ;
    END
  END w_mask_w1[315]
  PIN w_mask_w1[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.485 0.070 205.555 ;
    END
  END w_mask_w1[316]
  PIN w_mask_w1[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.045 0.070 206.115 ;
    END
  END w_mask_w1[317]
  PIN w_mask_w1[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.605 0.070 206.675 ;
    END
  END w_mask_w1[318]
  PIN w_mask_w1[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.165 0.070 207.235 ;
    END
  END w_mask_w1[319]
  PIN w_mask_w1[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.725 0.070 207.795 ;
    END
  END w_mask_w1[320]
  PIN w_mask_w1[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.285 0.070 208.355 ;
    END
  END w_mask_w1[321]
  PIN w_mask_w1[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.845 0.070 208.915 ;
    END
  END w_mask_w1[322]
  PIN w_mask_w1[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.405 0.070 209.475 ;
    END
  END w_mask_w1[323]
  PIN w_mask_w1[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.965 0.070 210.035 ;
    END
  END w_mask_w1[324]
  PIN w_mask_w1[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.525 0.070 210.595 ;
    END
  END w_mask_w1[325]
  PIN w_mask_w1[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.085 0.070 211.155 ;
    END
  END w_mask_w1[326]
  PIN w_mask_w1[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.645 0.070 211.715 ;
    END
  END w_mask_w1[327]
  PIN w_mask_w1[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.205 0.070 212.275 ;
    END
  END w_mask_w1[328]
  PIN w_mask_w1[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.765 0.070 212.835 ;
    END
  END w_mask_w1[329]
  PIN w_mask_w1[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.325 0.070 213.395 ;
    END
  END w_mask_w1[330]
  PIN w_mask_w1[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.885 0.070 213.955 ;
    END
  END w_mask_w1[331]
  PIN w_mask_w1[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.445 0.070 214.515 ;
    END
  END w_mask_w1[332]
  PIN w_mask_w1[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.005 0.070 215.075 ;
    END
  END w_mask_w1[333]
  PIN w_mask_w1[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.565 0.070 215.635 ;
    END
  END w_mask_w1[334]
  PIN w_mask_w1[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.125 0.070 216.195 ;
    END
  END w_mask_w1[335]
  PIN w_mask_w1[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.685 0.070 216.755 ;
    END
  END w_mask_w1[336]
  PIN w_mask_w1[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.245 0.070 217.315 ;
    END
  END w_mask_w1[337]
  PIN w_mask_w1[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.805 0.070 217.875 ;
    END
  END w_mask_w1[338]
  PIN w_mask_w1[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.365 0.070 218.435 ;
    END
  END w_mask_w1[339]
  PIN w_mask_w1[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.925 0.070 218.995 ;
    END
  END w_mask_w1[340]
  PIN w_mask_w1[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.485 0.070 219.555 ;
    END
  END w_mask_w1[341]
  PIN w_mask_w1[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.045 0.070 220.115 ;
    END
  END w_mask_w1[342]
  PIN w_mask_w1[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.605 0.070 220.675 ;
    END
  END w_mask_w1[343]
  PIN w_mask_w1[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.165 0.070 221.235 ;
    END
  END w_mask_w1[344]
  PIN w_mask_w1[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.725 0.070 221.795 ;
    END
  END w_mask_w1[345]
  PIN w_mask_w1[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.285 0.070 222.355 ;
    END
  END w_mask_w1[346]
  PIN w_mask_w1[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.845 0.070 222.915 ;
    END
  END w_mask_w1[347]
  PIN w_mask_w1[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.405 0.070 223.475 ;
    END
  END w_mask_w1[348]
  PIN w_mask_w1[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.965 0.070 224.035 ;
    END
  END w_mask_w1[349]
  PIN w_mask_w1[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.525 0.070 224.595 ;
    END
  END w_mask_w1[350]
  PIN w_mask_w1[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.085 0.070 225.155 ;
    END
  END w_mask_w1[351]
  PIN w_mask_w1[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.645 0.070 225.715 ;
    END
  END w_mask_w1[352]
  PIN w_mask_w1[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.205 0.070 226.275 ;
    END
  END w_mask_w1[353]
  PIN w_mask_w1[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.765 0.070 226.835 ;
    END
  END w_mask_w1[354]
  PIN w_mask_w1[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.325 0.070 227.395 ;
    END
  END w_mask_w1[355]
  PIN w_mask_w1[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.885 0.070 227.955 ;
    END
  END w_mask_w1[356]
  PIN w_mask_w1[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.445 0.070 228.515 ;
    END
  END w_mask_w1[357]
  PIN w_mask_w1[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.005 0.070 229.075 ;
    END
  END w_mask_w1[358]
  PIN w_mask_w1[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.565 0.070 229.635 ;
    END
  END w_mask_w1[359]
  PIN w_mask_w1[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.125 0.070 230.195 ;
    END
  END w_mask_w1[360]
  PIN w_mask_w1[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.685 0.070 230.755 ;
    END
  END w_mask_w1[361]
  PIN w_mask_w1[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.245 0.070 231.315 ;
    END
  END w_mask_w1[362]
  PIN w_mask_w1[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.805 0.070 231.875 ;
    END
  END w_mask_w1[363]
  PIN w_mask_w1[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.365 0.070 232.435 ;
    END
  END w_mask_w1[364]
  PIN w_mask_w1[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.925 0.070 232.995 ;
    END
  END w_mask_w1[365]
  PIN w_mask_w1[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.485 0.070 233.555 ;
    END
  END w_mask_w1[366]
  PIN w_mask_w1[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.045 0.070 234.115 ;
    END
  END w_mask_w1[367]
  PIN w_mask_w1[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.605 0.070 234.675 ;
    END
  END w_mask_w1[368]
  PIN w_mask_w1[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.165 0.070 235.235 ;
    END
  END w_mask_w1[369]
  PIN w_mask_w1[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.725 0.070 235.795 ;
    END
  END w_mask_w1[370]
  PIN w_mask_w1[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.285 0.070 236.355 ;
    END
  END w_mask_w1[371]
  PIN w_mask_w1[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.845 0.070 236.915 ;
    END
  END w_mask_w1[372]
  PIN w_mask_w1[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.405 0.070 237.475 ;
    END
  END w_mask_w1[373]
  PIN w_mask_w1[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.965 0.070 238.035 ;
    END
  END w_mask_w1[374]
  PIN w_mask_w1[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.525 0.070 238.595 ;
    END
  END w_mask_w1[375]
  PIN w_mask_w1[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.085 0.070 239.155 ;
    END
  END w_mask_w1[376]
  PIN w_mask_w1[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.645 0.070 239.715 ;
    END
  END w_mask_w1[377]
  PIN w_mask_w1[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.205 0.070 240.275 ;
    END
  END w_mask_w1[378]
  PIN w_mask_w1[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.765 0.070 240.835 ;
    END
  END w_mask_w1[379]
  PIN w_mask_w1[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.325 0.070 241.395 ;
    END
  END w_mask_w1[380]
  PIN w_mask_w1[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.885 0.070 241.955 ;
    END
  END w_mask_w1[381]
  PIN w_mask_w1[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.445 0.070 242.515 ;
    END
  END w_mask_w1[382]
  PIN w_mask_w1[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.005 0.070 243.075 ;
    END
  END w_mask_w1[383]
  PIN w_mask_w1[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.565 0.070 243.635 ;
    END
  END w_mask_w1[384]
  PIN w_mask_w1[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.125 0.070 244.195 ;
    END
  END w_mask_w1[385]
  PIN w_mask_w1[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.685 0.070 244.755 ;
    END
  END w_mask_w1[386]
  PIN w_mask_w1[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 245.245 0.070 245.315 ;
    END
  END w_mask_w1[387]
  PIN w_mask_w1[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 245.805 0.070 245.875 ;
    END
  END w_mask_w1[388]
  PIN w_mask_w1[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.365 0.070 246.435 ;
    END
  END w_mask_w1[389]
  PIN w_mask_w1[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.925 0.070 246.995 ;
    END
  END w_mask_w1[390]
  PIN w_mask_w1[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.485 0.070 247.555 ;
    END
  END w_mask_w1[391]
  PIN w_mask_w1[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.045 0.070 248.115 ;
    END
  END w_mask_w1[392]
  PIN w_mask_w1[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.605 0.070 248.675 ;
    END
  END w_mask_w1[393]
  PIN w_mask_w1[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.165 0.070 249.235 ;
    END
  END w_mask_w1[394]
  PIN w_mask_w1[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.725 0.070 249.795 ;
    END
  END w_mask_w1[395]
  PIN w_mask_w1[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.285 0.070 250.355 ;
    END
  END w_mask_w1[396]
  PIN w_mask_w1[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.845 0.070 250.915 ;
    END
  END w_mask_w1[397]
  PIN w_mask_w1[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.405 0.070 251.475 ;
    END
  END w_mask_w1[398]
  PIN w_mask_w1[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.965 0.070 252.035 ;
    END
  END w_mask_w1[399]
  PIN w_mask_w1[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.525 0.070 252.595 ;
    END
  END w_mask_w1[400]
  PIN w_mask_w1[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.085 0.070 253.155 ;
    END
  END w_mask_w1[401]
  PIN w_mask_w1[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.645 0.070 253.715 ;
    END
  END w_mask_w1[402]
  PIN w_mask_w1[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.205 0.070 254.275 ;
    END
  END w_mask_w1[403]
  PIN w_mask_w1[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.765 0.070 254.835 ;
    END
  END w_mask_w1[404]
  PIN w_mask_w1[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.325 0.070 255.395 ;
    END
  END w_mask_w1[405]
  PIN w_mask_w1[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.885 0.070 255.955 ;
    END
  END w_mask_w1[406]
  PIN w_mask_w1[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.445 0.070 256.515 ;
    END
  END w_mask_w1[407]
  PIN w_mask_w1[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.005 0.070 257.075 ;
    END
  END w_mask_w1[408]
  PIN w_mask_w1[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.565 0.070 257.635 ;
    END
  END w_mask_w1[409]
  PIN w_mask_w1[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.125 0.070 258.195 ;
    END
  END w_mask_w1[410]
  PIN w_mask_w1[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.685 0.070 258.755 ;
    END
  END w_mask_w1[411]
  PIN w_mask_w1[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.245 0.070 259.315 ;
    END
  END w_mask_w1[412]
  PIN w_mask_w1[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.805 0.070 259.875 ;
    END
  END w_mask_w1[413]
  PIN w_mask_w1[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.365 0.070 260.435 ;
    END
  END w_mask_w1[414]
  PIN w_mask_w1[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.925 0.070 260.995 ;
    END
  END w_mask_w1[415]
  PIN w_mask_w1[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 261.485 0.070 261.555 ;
    END
  END w_mask_w1[416]
  PIN w_mask_w1[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.045 0.070 262.115 ;
    END
  END w_mask_w1[417]
  PIN w_mask_w1[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.605 0.070 262.675 ;
    END
  END w_mask_w1[418]
  PIN w_mask_w1[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.165 0.070 263.235 ;
    END
  END w_mask_w1[419]
  PIN w_mask_w1[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.725 0.070 263.795 ;
    END
  END w_mask_w1[420]
  PIN w_mask_w1[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.285 0.070 264.355 ;
    END
  END w_mask_w1[421]
  PIN w_mask_w1[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.845 0.070 264.915 ;
    END
  END w_mask_w1[422]
  PIN w_mask_w1[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 265.405 0.070 265.475 ;
    END
  END w_mask_w1[423]
  PIN w_mask_w1[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 265.965 0.070 266.035 ;
    END
  END w_mask_w1[424]
  PIN w_mask_w1[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.525 0.070 266.595 ;
    END
  END w_mask_w1[425]
  PIN w_mask_w1[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.085 0.070 267.155 ;
    END
  END w_mask_w1[426]
  PIN w_mask_w1[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.645 0.070 267.715 ;
    END
  END w_mask_w1[427]
  PIN w_mask_w1[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.205 0.070 268.275 ;
    END
  END w_mask_w1[428]
  PIN w_mask_w1[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.765 0.070 268.835 ;
    END
  END w_mask_w1[429]
  PIN w_mask_w1[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.325 0.070 269.395 ;
    END
  END w_mask_w1[430]
  PIN w_mask_w1[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.885 0.070 269.955 ;
    END
  END w_mask_w1[431]
  PIN w_mask_w1[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.445 0.070 270.515 ;
    END
  END w_mask_w1[432]
  PIN w_mask_w1[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.005 0.070 271.075 ;
    END
  END w_mask_w1[433]
  PIN w_mask_w1[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.565 0.070 271.635 ;
    END
  END w_mask_w1[434]
  PIN w_mask_w1[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.125 0.070 272.195 ;
    END
  END w_mask_w1[435]
  PIN w_mask_w1[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.685 0.070 272.755 ;
    END
  END w_mask_w1[436]
  PIN w_mask_w1[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.245 0.070 273.315 ;
    END
  END w_mask_w1[437]
  PIN w_mask_w1[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.805 0.070 273.875 ;
    END
  END w_mask_w1[438]
  PIN w_mask_w1[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.365 0.070 274.435 ;
    END
  END w_mask_w1[439]
  PIN w_mask_w1[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.925 0.070 274.995 ;
    END
  END w_mask_w1[440]
  PIN w_mask_w1[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.485 0.070 275.555 ;
    END
  END w_mask_w1[441]
  PIN w_mask_w1[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.045 0.070 276.115 ;
    END
  END w_mask_w1[442]
  PIN w_mask_w1[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.605 0.070 276.675 ;
    END
  END w_mask_w1[443]
  PIN w_mask_w1[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.165 0.070 277.235 ;
    END
  END w_mask_w1[444]
  PIN w_mask_w1[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.725 0.070 277.795 ;
    END
  END w_mask_w1[445]
  PIN w_mask_w1[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.285 0.070 278.355 ;
    END
  END w_mask_w1[446]
  PIN w_mask_w1[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.845 0.070 278.915 ;
    END
  END w_mask_w1[447]
  PIN w_mask_w1[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.405 0.070 279.475 ;
    END
  END w_mask_w1[448]
  PIN w_mask_w1[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.965 0.070 280.035 ;
    END
  END w_mask_w1[449]
  PIN w_mask_w1[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.525 0.070 280.595 ;
    END
  END w_mask_w1[450]
  PIN w_mask_w1[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.085 0.070 281.155 ;
    END
  END w_mask_w1[451]
  PIN w_mask_w1[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.645 0.070 281.715 ;
    END
  END w_mask_w1[452]
  PIN w_mask_w1[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.205 0.070 282.275 ;
    END
  END w_mask_w1[453]
  PIN w_mask_w1[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.765 0.070 282.835 ;
    END
  END w_mask_w1[454]
  PIN w_mask_w1[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.325 0.070 283.395 ;
    END
  END w_mask_w1[455]
  PIN w_mask_w1[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.885 0.070 283.955 ;
    END
  END w_mask_w1[456]
  PIN w_mask_w1[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.445 0.070 284.515 ;
    END
  END w_mask_w1[457]
  PIN w_mask_w1[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.005 0.070 285.075 ;
    END
  END w_mask_w1[458]
  PIN w_mask_w1[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.565 0.070 285.635 ;
    END
  END w_mask_w1[459]
  PIN w_mask_w1[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.125 0.070 286.195 ;
    END
  END w_mask_w1[460]
  PIN w_mask_w1[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.685 0.070 286.755 ;
    END
  END w_mask_w1[461]
  PIN w_mask_w1[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.245 0.070 287.315 ;
    END
  END w_mask_w1[462]
  PIN w_mask_w1[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.805 0.070 287.875 ;
    END
  END w_mask_w1[463]
  PIN w_mask_w1[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.365 0.070 288.435 ;
    END
  END w_mask_w1[464]
  PIN w_mask_w1[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.925 0.070 288.995 ;
    END
  END w_mask_w1[465]
  PIN w_mask_w1[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.485 0.070 289.555 ;
    END
  END w_mask_w1[466]
  PIN w_mask_w1[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.045 0.070 290.115 ;
    END
  END w_mask_w1[467]
  PIN w_mask_w1[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.605 0.070 290.675 ;
    END
  END w_mask_w1[468]
  PIN w_mask_w1[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.165 0.070 291.235 ;
    END
  END w_mask_w1[469]
  PIN w_mask_w1[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.725 0.070 291.795 ;
    END
  END w_mask_w1[470]
  PIN w_mask_w1[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.285 0.070 292.355 ;
    END
  END w_mask_w1[471]
  PIN w_mask_w1[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.845 0.070 292.915 ;
    END
  END w_mask_w1[472]
  PIN w_mask_w1[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.405 0.070 293.475 ;
    END
  END w_mask_w1[473]
  PIN w_mask_w1[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.965 0.070 294.035 ;
    END
  END w_mask_w1[474]
  PIN w_mask_w1[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.525 0.070 294.595 ;
    END
  END w_mask_w1[475]
  PIN w_mask_w1[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.085 0.070 295.155 ;
    END
  END w_mask_w1[476]
  PIN w_mask_w1[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.645 0.070 295.715 ;
    END
  END w_mask_w1[477]
  PIN w_mask_w1[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.205 0.070 296.275 ;
    END
  END w_mask_w1[478]
  PIN w_mask_w1[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.765 0.070 296.835 ;
    END
  END w_mask_w1[479]
  PIN w_mask_w1[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.325 0.070 297.395 ;
    END
  END w_mask_w1[480]
  PIN w_mask_w1[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.885 0.070 297.955 ;
    END
  END w_mask_w1[481]
  PIN w_mask_w1[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.445 0.070 298.515 ;
    END
  END w_mask_w1[482]
  PIN w_mask_w1[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.005 0.070 299.075 ;
    END
  END w_mask_w1[483]
  PIN w_mask_w1[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.565 0.070 299.635 ;
    END
  END w_mask_w1[484]
  PIN w_mask_w1[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.125 0.070 300.195 ;
    END
  END w_mask_w1[485]
  PIN w_mask_w1[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.685 0.070 300.755 ;
    END
  END w_mask_w1[486]
  PIN w_mask_w1[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.245 0.070 301.315 ;
    END
  END w_mask_w1[487]
  PIN w_mask_w1[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.805 0.070 301.875 ;
    END
  END w_mask_w1[488]
  PIN w_mask_w1[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.365 0.070 302.435 ;
    END
  END w_mask_w1[489]
  PIN w_mask_w1[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.925 0.070 302.995 ;
    END
  END w_mask_w1[490]
  PIN w_mask_w1[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.485 0.070 303.555 ;
    END
  END w_mask_w1[491]
  PIN w_mask_w1[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.045 0.070 304.115 ;
    END
  END w_mask_w1[492]
  PIN w_mask_w1[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.605 0.070 304.675 ;
    END
  END w_mask_w1[493]
  PIN w_mask_w1[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.165 0.070 305.235 ;
    END
  END w_mask_w1[494]
  PIN w_mask_w1[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.725 0.070 305.795 ;
    END
  END w_mask_w1[495]
  PIN w_mask_w1[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.285 0.070 306.355 ;
    END
  END w_mask_w1[496]
  PIN w_mask_w1[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.845 0.070 306.915 ;
    END
  END w_mask_w1[497]
  PIN w_mask_w1[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.405 0.070 307.475 ;
    END
  END w_mask_w1[498]
  PIN w_mask_w1[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.965 0.070 308.035 ;
    END
  END w_mask_w1[499]
  PIN w_mask_w1[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.525 0.070 308.595 ;
    END
  END w_mask_w1[500]
  PIN w_mask_w1[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.085 0.070 309.155 ;
    END
  END w_mask_w1[501]
  PIN w_mask_w1[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.645 0.070 309.715 ;
    END
  END w_mask_w1[502]
  PIN w_mask_w1[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.205 0.070 310.275 ;
    END
  END w_mask_w1[503]
  PIN w_mask_w1[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.765 0.070 310.835 ;
    END
  END w_mask_w1[504]
  PIN w_mask_w1[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.325 0.070 311.395 ;
    END
  END w_mask_w1[505]
  PIN w_mask_w1[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.885 0.070 311.955 ;
    END
  END w_mask_w1[506]
  PIN w_mask_w1[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.445 0.070 312.515 ;
    END
  END w_mask_w1[507]
  PIN w_mask_w1[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.005 0.070 313.075 ;
    END
  END w_mask_w1[508]
  PIN w_mask_w1[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.565 0.070 313.635 ;
    END
  END w_mask_w1[509]
  PIN w_mask_w1[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.125 0.070 314.195 ;
    END
  END w_mask_w1[510]
  PIN w_mask_w1[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.685 0.070 314.755 ;
    END
  END w_mask_w1[511]
  PIN rd_out_r1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.405 0.070 342.475 ;
    END
  END rd_out_r1[0]
  PIN rd_out_r1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.965 0.070 343.035 ;
    END
  END rd_out_r1[1]
  PIN rd_out_r1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.525 0.070 343.595 ;
    END
  END rd_out_r1[2]
  PIN rd_out_r1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.085 0.070 344.155 ;
    END
  END rd_out_r1[3]
  PIN rd_out_r1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.645 0.070 344.715 ;
    END
  END rd_out_r1[4]
  PIN rd_out_r1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.205 0.070 345.275 ;
    END
  END rd_out_r1[5]
  PIN rd_out_r1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.765 0.070 345.835 ;
    END
  END rd_out_r1[6]
  PIN rd_out_r1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.325 0.070 346.395 ;
    END
  END rd_out_r1[7]
  PIN rd_out_r1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.885 0.070 346.955 ;
    END
  END rd_out_r1[8]
  PIN rd_out_r1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.445 0.070 347.515 ;
    END
  END rd_out_r1[9]
  PIN rd_out_r1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.005 0.070 348.075 ;
    END
  END rd_out_r1[10]
  PIN rd_out_r1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.565 0.070 348.635 ;
    END
  END rd_out_r1[11]
  PIN rd_out_r1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.125 0.070 349.195 ;
    END
  END rd_out_r1[12]
  PIN rd_out_r1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.685 0.070 349.755 ;
    END
  END rd_out_r1[13]
  PIN rd_out_r1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.245 0.070 350.315 ;
    END
  END rd_out_r1[14]
  PIN rd_out_r1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.805 0.070 350.875 ;
    END
  END rd_out_r1[15]
  PIN rd_out_r1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.365 0.070 351.435 ;
    END
  END rd_out_r1[16]
  PIN rd_out_r1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.925 0.070 351.995 ;
    END
  END rd_out_r1[17]
  PIN rd_out_r1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.485 0.070 352.555 ;
    END
  END rd_out_r1[18]
  PIN rd_out_r1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.045 0.070 353.115 ;
    END
  END rd_out_r1[19]
  PIN rd_out_r1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.605 0.070 353.675 ;
    END
  END rd_out_r1[20]
  PIN rd_out_r1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.165 0.070 354.235 ;
    END
  END rd_out_r1[21]
  PIN rd_out_r1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.725 0.070 354.795 ;
    END
  END rd_out_r1[22]
  PIN rd_out_r1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.285 0.070 355.355 ;
    END
  END rd_out_r1[23]
  PIN rd_out_r1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.845 0.070 355.915 ;
    END
  END rd_out_r1[24]
  PIN rd_out_r1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.405 0.070 356.475 ;
    END
  END rd_out_r1[25]
  PIN rd_out_r1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.965 0.070 357.035 ;
    END
  END rd_out_r1[26]
  PIN rd_out_r1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.525 0.070 357.595 ;
    END
  END rd_out_r1[27]
  PIN rd_out_r1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.085 0.070 358.155 ;
    END
  END rd_out_r1[28]
  PIN rd_out_r1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.645 0.070 358.715 ;
    END
  END rd_out_r1[29]
  PIN rd_out_r1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.205 0.070 359.275 ;
    END
  END rd_out_r1[30]
  PIN rd_out_r1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.765 0.070 359.835 ;
    END
  END rd_out_r1[31]
  PIN rd_out_r1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.325 0.070 360.395 ;
    END
  END rd_out_r1[32]
  PIN rd_out_r1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.885 0.070 360.955 ;
    END
  END rd_out_r1[33]
  PIN rd_out_r1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 361.445 0.070 361.515 ;
    END
  END rd_out_r1[34]
  PIN rd_out_r1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.005 0.070 362.075 ;
    END
  END rd_out_r1[35]
  PIN rd_out_r1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.565 0.070 362.635 ;
    END
  END rd_out_r1[36]
  PIN rd_out_r1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.125 0.070 363.195 ;
    END
  END rd_out_r1[37]
  PIN rd_out_r1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.685 0.070 363.755 ;
    END
  END rd_out_r1[38]
  PIN rd_out_r1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.245 0.070 364.315 ;
    END
  END rd_out_r1[39]
  PIN rd_out_r1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.805 0.070 364.875 ;
    END
  END rd_out_r1[40]
  PIN rd_out_r1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.365 0.070 365.435 ;
    END
  END rd_out_r1[41]
  PIN rd_out_r1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.925 0.070 365.995 ;
    END
  END rd_out_r1[42]
  PIN rd_out_r1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 366.485 0.070 366.555 ;
    END
  END rd_out_r1[43]
  PIN rd_out_r1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.045 0.070 367.115 ;
    END
  END rd_out_r1[44]
  PIN rd_out_r1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.605 0.070 367.675 ;
    END
  END rd_out_r1[45]
  PIN rd_out_r1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.165 0.070 368.235 ;
    END
  END rd_out_r1[46]
  PIN rd_out_r1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.725 0.070 368.795 ;
    END
  END rd_out_r1[47]
  PIN rd_out_r1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.285 0.070 369.355 ;
    END
  END rd_out_r1[48]
  PIN rd_out_r1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.845 0.070 369.915 ;
    END
  END rd_out_r1[49]
  PIN rd_out_r1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.405 0.070 370.475 ;
    END
  END rd_out_r1[50]
  PIN rd_out_r1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.965 0.070 371.035 ;
    END
  END rd_out_r1[51]
  PIN rd_out_r1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 371.525 0.070 371.595 ;
    END
  END rd_out_r1[52]
  PIN rd_out_r1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.085 0.070 372.155 ;
    END
  END rd_out_r1[53]
  PIN rd_out_r1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.645 0.070 372.715 ;
    END
  END rd_out_r1[54]
  PIN rd_out_r1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.205 0.070 373.275 ;
    END
  END rd_out_r1[55]
  PIN rd_out_r1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.765 0.070 373.835 ;
    END
  END rd_out_r1[56]
  PIN rd_out_r1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.325 0.070 374.395 ;
    END
  END rd_out_r1[57]
  PIN rd_out_r1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.885 0.070 374.955 ;
    END
  END rd_out_r1[58]
  PIN rd_out_r1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 375.445 0.070 375.515 ;
    END
  END rd_out_r1[59]
  PIN rd_out_r1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.005 0.070 376.075 ;
    END
  END rd_out_r1[60]
  PIN rd_out_r1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.565 0.070 376.635 ;
    END
  END rd_out_r1[61]
  PIN rd_out_r1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.125 0.070 377.195 ;
    END
  END rd_out_r1[62]
  PIN rd_out_r1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.685 0.070 377.755 ;
    END
  END rd_out_r1[63]
  PIN rd_out_r1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.245 0.070 378.315 ;
    END
  END rd_out_r1[64]
  PIN rd_out_r1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.805 0.070 378.875 ;
    END
  END rd_out_r1[65]
  PIN rd_out_r1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.365 0.070 379.435 ;
    END
  END rd_out_r1[66]
  PIN rd_out_r1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.925 0.070 379.995 ;
    END
  END rd_out_r1[67]
  PIN rd_out_r1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 380.485 0.070 380.555 ;
    END
  END rd_out_r1[68]
  PIN rd_out_r1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.045 0.070 381.115 ;
    END
  END rd_out_r1[69]
  PIN rd_out_r1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.605 0.070 381.675 ;
    END
  END rd_out_r1[70]
  PIN rd_out_r1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 382.165 0.070 382.235 ;
    END
  END rd_out_r1[71]
  PIN rd_out_r1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 382.725 0.070 382.795 ;
    END
  END rd_out_r1[72]
  PIN rd_out_r1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.285 0.070 383.355 ;
    END
  END rd_out_r1[73]
  PIN rd_out_r1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.845 0.070 383.915 ;
    END
  END rd_out_r1[74]
  PIN rd_out_r1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.405 0.070 384.475 ;
    END
  END rd_out_r1[75]
  PIN rd_out_r1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.965 0.070 385.035 ;
    END
  END rd_out_r1[76]
  PIN rd_out_r1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.525 0.070 385.595 ;
    END
  END rd_out_r1[77]
  PIN rd_out_r1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.085 0.070 386.155 ;
    END
  END rd_out_r1[78]
  PIN rd_out_r1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.645 0.070 386.715 ;
    END
  END rd_out_r1[79]
  PIN rd_out_r1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.205 0.070 387.275 ;
    END
  END rd_out_r1[80]
  PIN rd_out_r1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.765 0.070 387.835 ;
    END
  END rd_out_r1[81]
  PIN rd_out_r1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.325 0.070 388.395 ;
    END
  END rd_out_r1[82]
  PIN rd_out_r1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.885 0.070 388.955 ;
    END
  END rd_out_r1[83]
  PIN rd_out_r1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 389.445 0.070 389.515 ;
    END
  END rd_out_r1[84]
  PIN rd_out_r1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.005 0.070 390.075 ;
    END
  END rd_out_r1[85]
  PIN rd_out_r1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.565 0.070 390.635 ;
    END
  END rd_out_r1[86]
  PIN rd_out_r1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.125 0.070 391.195 ;
    END
  END rd_out_r1[87]
  PIN rd_out_r1[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.685 0.070 391.755 ;
    END
  END rd_out_r1[88]
  PIN rd_out_r1[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.245 0.070 392.315 ;
    END
  END rd_out_r1[89]
  PIN rd_out_r1[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.805 0.070 392.875 ;
    END
  END rd_out_r1[90]
  PIN rd_out_r1[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.365 0.070 393.435 ;
    END
  END rd_out_r1[91]
  PIN rd_out_r1[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.925 0.070 393.995 ;
    END
  END rd_out_r1[92]
  PIN rd_out_r1[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.485 0.070 394.555 ;
    END
  END rd_out_r1[93]
  PIN rd_out_r1[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.045 0.070 395.115 ;
    END
  END rd_out_r1[94]
  PIN rd_out_r1[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.605 0.070 395.675 ;
    END
  END rd_out_r1[95]
  PIN rd_out_r1[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.165 0.070 396.235 ;
    END
  END rd_out_r1[96]
  PIN rd_out_r1[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.725 0.070 396.795 ;
    END
  END rd_out_r1[97]
  PIN rd_out_r1[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.285 0.070 397.355 ;
    END
  END rd_out_r1[98]
  PIN rd_out_r1[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.845 0.070 397.915 ;
    END
  END rd_out_r1[99]
  PIN rd_out_r1[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.405 0.070 398.475 ;
    END
  END rd_out_r1[100]
  PIN rd_out_r1[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.965 0.070 399.035 ;
    END
  END rd_out_r1[101]
  PIN rd_out_r1[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.525 0.070 399.595 ;
    END
  END rd_out_r1[102]
  PIN rd_out_r1[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 400.085 0.070 400.155 ;
    END
  END rd_out_r1[103]
  PIN rd_out_r1[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 400.645 0.070 400.715 ;
    END
  END rd_out_r1[104]
  PIN rd_out_r1[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 401.205 0.070 401.275 ;
    END
  END rd_out_r1[105]
  PIN rd_out_r1[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 401.765 0.070 401.835 ;
    END
  END rd_out_r1[106]
  PIN rd_out_r1[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 402.325 0.070 402.395 ;
    END
  END rd_out_r1[107]
  PIN rd_out_r1[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 402.885 0.070 402.955 ;
    END
  END rd_out_r1[108]
  PIN rd_out_r1[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 403.445 0.070 403.515 ;
    END
  END rd_out_r1[109]
  PIN rd_out_r1[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 404.005 0.070 404.075 ;
    END
  END rd_out_r1[110]
  PIN rd_out_r1[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 404.565 0.070 404.635 ;
    END
  END rd_out_r1[111]
  PIN rd_out_r1[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 405.125 0.070 405.195 ;
    END
  END rd_out_r1[112]
  PIN rd_out_r1[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 405.685 0.070 405.755 ;
    END
  END rd_out_r1[113]
  PIN rd_out_r1[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 406.245 0.070 406.315 ;
    END
  END rd_out_r1[114]
  PIN rd_out_r1[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 406.805 0.070 406.875 ;
    END
  END rd_out_r1[115]
  PIN rd_out_r1[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 407.365 0.070 407.435 ;
    END
  END rd_out_r1[116]
  PIN rd_out_r1[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 407.925 0.070 407.995 ;
    END
  END rd_out_r1[117]
  PIN rd_out_r1[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 408.485 0.070 408.555 ;
    END
  END rd_out_r1[118]
  PIN rd_out_r1[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 409.045 0.070 409.115 ;
    END
  END rd_out_r1[119]
  PIN rd_out_r1[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 409.605 0.070 409.675 ;
    END
  END rd_out_r1[120]
  PIN rd_out_r1[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 410.165 0.070 410.235 ;
    END
  END rd_out_r1[121]
  PIN rd_out_r1[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 410.725 0.070 410.795 ;
    END
  END rd_out_r1[122]
  PIN rd_out_r1[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 411.285 0.070 411.355 ;
    END
  END rd_out_r1[123]
  PIN rd_out_r1[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 411.845 0.070 411.915 ;
    END
  END rd_out_r1[124]
  PIN rd_out_r1[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 412.405 0.070 412.475 ;
    END
  END rd_out_r1[125]
  PIN rd_out_r1[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 412.965 0.070 413.035 ;
    END
  END rd_out_r1[126]
  PIN rd_out_r1[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 413.525 0.070 413.595 ;
    END
  END rd_out_r1[127]
  PIN rd_out_r1[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 414.085 0.070 414.155 ;
    END
  END rd_out_r1[128]
  PIN rd_out_r1[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 414.645 0.070 414.715 ;
    END
  END rd_out_r1[129]
  PIN rd_out_r1[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 415.205 0.070 415.275 ;
    END
  END rd_out_r1[130]
  PIN rd_out_r1[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 415.765 0.070 415.835 ;
    END
  END rd_out_r1[131]
  PIN rd_out_r1[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 416.325 0.070 416.395 ;
    END
  END rd_out_r1[132]
  PIN rd_out_r1[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 416.885 0.070 416.955 ;
    END
  END rd_out_r1[133]
  PIN rd_out_r1[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 417.445 0.070 417.515 ;
    END
  END rd_out_r1[134]
  PIN rd_out_r1[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 418.005 0.070 418.075 ;
    END
  END rd_out_r1[135]
  PIN rd_out_r1[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 418.565 0.070 418.635 ;
    END
  END rd_out_r1[136]
  PIN rd_out_r1[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 419.125 0.070 419.195 ;
    END
  END rd_out_r1[137]
  PIN rd_out_r1[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 419.685 0.070 419.755 ;
    END
  END rd_out_r1[138]
  PIN rd_out_r1[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 420.245 0.070 420.315 ;
    END
  END rd_out_r1[139]
  PIN rd_out_r1[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 420.805 0.070 420.875 ;
    END
  END rd_out_r1[140]
  PIN rd_out_r1[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 421.365 0.070 421.435 ;
    END
  END rd_out_r1[141]
  PIN rd_out_r1[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 421.925 0.070 421.995 ;
    END
  END rd_out_r1[142]
  PIN rd_out_r1[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 422.485 0.070 422.555 ;
    END
  END rd_out_r1[143]
  PIN rd_out_r1[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 423.045 0.070 423.115 ;
    END
  END rd_out_r1[144]
  PIN rd_out_r1[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 423.605 0.070 423.675 ;
    END
  END rd_out_r1[145]
  PIN rd_out_r1[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 424.165 0.070 424.235 ;
    END
  END rd_out_r1[146]
  PIN rd_out_r1[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 424.725 0.070 424.795 ;
    END
  END rd_out_r1[147]
  PIN rd_out_r1[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 425.285 0.070 425.355 ;
    END
  END rd_out_r1[148]
  PIN rd_out_r1[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 425.845 0.070 425.915 ;
    END
  END rd_out_r1[149]
  PIN rd_out_r1[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 426.405 0.070 426.475 ;
    END
  END rd_out_r1[150]
  PIN rd_out_r1[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 426.965 0.070 427.035 ;
    END
  END rd_out_r1[151]
  PIN rd_out_r1[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 427.525 0.070 427.595 ;
    END
  END rd_out_r1[152]
  PIN rd_out_r1[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 428.085 0.070 428.155 ;
    END
  END rd_out_r1[153]
  PIN rd_out_r1[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 428.645 0.070 428.715 ;
    END
  END rd_out_r1[154]
  PIN rd_out_r1[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 429.205 0.070 429.275 ;
    END
  END rd_out_r1[155]
  PIN rd_out_r1[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 429.765 0.070 429.835 ;
    END
  END rd_out_r1[156]
  PIN rd_out_r1[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 430.325 0.070 430.395 ;
    END
  END rd_out_r1[157]
  PIN rd_out_r1[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 430.885 0.070 430.955 ;
    END
  END rd_out_r1[158]
  PIN rd_out_r1[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 431.445 0.070 431.515 ;
    END
  END rd_out_r1[159]
  PIN rd_out_r1[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 432.005 0.070 432.075 ;
    END
  END rd_out_r1[160]
  PIN rd_out_r1[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 432.565 0.070 432.635 ;
    END
  END rd_out_r1[161]
  PIN rd_out_r1[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 433.125 0.070 433.195 ;
    END
  END rd_out_r1[162]
  PIN rd_out_r1[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 433.685 0.070 433.755 ;
    END
  END rd_out_r1[163]
  PIN rd_out_r1[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 434.245 0.070 434.315 ;
    END
  END rd_out_r1[164]
  PIN rd_out_r1[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 434.805 0.070 434.875 ;
    END
  END rd_out_r1[165]
  PIN rd_out_r1[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 435.365 0.070 435.435 ;
    END
  END rd_out_r1[166]
  PIN rd_out_r1[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 435.925 0.070 435.995 ;
    END
  END rd_out_r1[167]
  PIN rd_out_r1[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 436.485 0.070 436.555 ;
    END
  END rd_out_r1[168]
  PIN rd_out_r1[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 437.045 0.070 437.115 ;
    END
  END rd_out_r1[169]
  PIN rd_out_r1[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 437.605 0.070 437.675 ;
    END
  END rd_out_r1[170]
  PIN rd_out_r1[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 438.165 0.070 438.235 ;
    END
  END rd_out_r1[171]
  PIN rd_out_r1[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 438.725 0.070 438.795 ;
    END
  END rd_out_r1[172]
  PIN rd_out_r1[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 439.285 0.070 439.355 ;
    END
  END rd_out_r1[173]
  PIN rd_out_r1[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 439.845 0.070 439.915 ;
    END
  END rd_out_r1[174]
  PIN rd_out_r1[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 440.405 0.070 440.475 ;
    END
  END rd_out_r1[175]
  PIN rd_out_r1[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 440.965 0.070 441.035 ;
    END
  END rd_out_r1[176]
  PIN rd_out_r1[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 441.525 0.070 441.595 ;
    END
  END rd_out_r1[177]
  PIN rd_out_r1[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 442.085 0.070 442.155 ;
    END
  END rd_out_r1[178]
  PIN rd_out_r1[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 442.645 0.070 442.715 ;
    END
  END rd_out_r1[179]
  PIN rd_out_r1[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 443.205 0.070 443.275 ;
    END
  END rd_out_r1[180]
  PIN rd_out_r1[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 443.765 0.070 443.835 ;
    END
  END rd_out_r1[181]
  PIN rd_out_r1[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 444.325 0.070 444.395 ;
    END
  END rd_out_r1[182]
  PIN rd_out_r1[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 444.885 0.070 444.955 ;
    END
  END rd_out_r1[183]
  PIN rd_out_r1[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 445.445 0.070 445.515 ;
    END
  END rd_out_r1[184]
  PIN rd_out_r1[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 446.005 0.070 446.075 ;
    END
  END rd_out_r1[185]
  PIN rd_out_r1[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 446.565 0.070 446.635 ;
    END
  END rd_out_r1[186]
  PIN rd_out_r1[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 447.125 0.070 447.195 ;
    END
  END rd_out_r1[187]
  PIN rd_out_r1[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 447.685 0.070 447.755 ;
    END
  END rd_out_r1[188]
  PIN rd_out_r1[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 448.245 0.070 448.315 ;
    END
  END rd_out_r1[189]
  PIN rd_out_r1[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 448.805 0.070 448.875 ;
    END
  END rd_out_r1[190]
  PIN rd_out_r1[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 449.365 0.070 449.435 ;
    END
  END rd_out_r1[191]
  PIN rd_out_r1[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 449.925 0.070 449.995 ;
    END
  END rd_out_r1[192]
  PIN rd_out_r1[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 450.485 0.070 450.555 ;
    END
  END rd_out_r1[193]
  PIN rd_out_r1[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 451.045 0.070 451.115 ;
    END
  END rd_out_r1[194]
  PIN rd_out_r1[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 451.605 0.070 451.675 ;
    END
  END rd_out_r1[195]
  PIN rd_out_r1[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 452.165 0.070 452.235 ;
    END
  END rd_out_r1[196]
  PIN rd_out_r1[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 452.725 0.070 452.795 ;
    END
  END rd_out_r1[197]
  PIN rd_out_r1[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 453.285 0.070 453.355 ;
    END
  END rd_out_r1[198]
  PIN rd_out_r1[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 453.845 0.070 453.915 ;
    END
  END rd_out_r1[199]
  PIN rd_out_r1[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 454.405 0.070 454.475 ;
    END
  END rd_out_r1[200]
  PIN rd_out_r1[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 454.965 0.070 455.035 ;
    END
  END rd_out_r1[201]
  PIN rd_out_r1[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 455.525 0.070 455.595 ;
    END
  END rd_out_r1[202]
  PIN rd_out_r1[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 456.085 0.070 456.155 ;
    END
  END rd_out_r1[203]
  PIN rd_out_r1[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 456.645 0.070 456.715 ;
    END
  END rd_out_r1[204]
  PIN rd_out_r1[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 457.205 0.070 457.275 ;
    END
  END rd_out_r1[205]
  PIN rd_out_r1[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 457.765 0.070 457.835 ;
    END
  END rd_out_r1[206]
  PIN rd_out_r1[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 458.325 0.070 458.395 ;
    END
  END rd_out_r1[207]
  PIN rd_out_r1[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 458.885 0.070 458.955 ;
    END
  END rd_out_r1[208]
  PIN rd_out_r1[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 459.445 0.070 459.515 ;
    END
  END rd_out_r1[209]
  PIN rd_out_r1[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 460.005 0.070 460.075 ;
    END
  END rd_out_r1[210]
  PIN rd_out_r1[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 460.565 0.070 460.635 ;
    END
  END rd_out_r1[211]
  PIN rd_out_r1[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 461.125 0.070 461.195 ;
    END
  END rd_out_r1[212]
  PIN rd_out_r1[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 461.685 0.070 461.755 ;
    END
  END rd_out_r1[213]
  PIN rd_out_r1[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 462.245 0.070 462.315 ;
    END
  END rd_out_r1[214]
  PIN rd_out_r1[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 462.805 0.070 462.875 ;
    END
  END rd_out_r1[215]
  PIN rd_out_r1[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 463.365 0.070 463.435 ;
    END
  END rd_out_r1[216]
  PIN rd_out_r1[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 463.925 0.070 463.995 ;
    END
  END rd_out_r1[217]
  PIN rd_out_r1[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 464.485 0.070 464.555 ;
    END
  END rd_out_r1[218]
  PIN rd_out_r1[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 465.045 0.070 465.115 ;
    END
  END rd_out_r1[219]
  PIN rd_out_r1[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 465.605 0.070 465.675 ;
    END
  END rd_out_r1[220]
  PIN rd_out_r1[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 466.165 0.070 466.235 ;
    END
  END rd_out_r1[221]
  PIN rd_out_r1[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 466.725 0.070 466.795 ;
    END
  END rd_out_r1[222]
  PIN rd_out_r1[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 467.285 0.070 467.355 ;
    END
  END rd_out_r1[223]
  PIN rd_out_r1[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 467.845 0.070 467.915 ;
    END
  END rd_out_r1[224]
  PIN rd_out_r1[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 468.405 0.070 468.475 ;
    END
  END rd_out_r1[225]
  PIN rd_out_r1[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 468.965 0.070 469.035 ;
    END
  END rd_out_r1[226]
  PIN rd_out_r1[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 469.525 0.070 469.595 ;
    END
  END rd_out_r1[227]
  PIN rd_out_r1[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 470.085 0.070 470.155 ;
    END
  END rd_out_r1[228]
  PIN rd_out_r1[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 470.645 0.070 470.715 ;
    END
  END rd_out_r1[229]
  PIN rd_out_r1[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 471.205 0.070 471.275 ;
    END
  END rd_out_r1[230]
  PIN rd_out_r1[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 471.765 0.070 471.835 ;
    END
  END rd_out_r1[231]
  PIN rd_out_r1[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 472.325 0.070 472.395 ;
    END
  END rd_out_r1[232]
  PIN rd_out_r1[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 472.885 0.070 472.955 ;
    END
  END rd_out_r1[233]
  PIN rd_out_r1[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 473.445 0.070 473.515 ;
    END
  END rd_out_r1[234]
  PIN rd_out_r1[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 474.005 0.070 474.075 ;
    END
  END rd_out_r1[235]
  PIN rd_out_r1[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 474.565 0.070 474.635 ;
    END
  END rd_out_r1[236]
  PIN rd_out_r1[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 475.125 0.070 475.195 ;
    END
  END rd_out_r1[237]
  PIN rd_out_r1[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 475.685 0.070 475.755 ;
    END
  END rd_out_r1[238]
  PIN rd_out_r1[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 476.245 0.070 476.315 ;
    END
  END rd_out_r1[239]
  PIN rd_out_r1[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 476.805 0.070 476.875 ;
    END
  END rd_out_r1[240]
  PIN rd_out_r1[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 477.365 0.070 477.435 ;
    END
  END rd_out_r1[241]
  PIN rd_out_r1[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 477.925 0.070 477.995 ;
    END
  END rd_out_r1[242]
  PIN rd_out_r1[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 478.485 0.070 478.555 ;
    END
  END rd_out_r1[243]
  PIN rd_out_r1[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 479.045 0.070 479.115 ;
    END
  END rd_out_r1[244]
  PIN rd_out_r1[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 479.605 0.070 479.675 ;
    END
  END rd_out_r1[245]
  PIN rd_out_r1[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 480.165 0.070 480.235 ;
    END
  END rd_out_r1[246]
  PIN rd_out_r1[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 480.725 0.070 480.795 ;
    END
  END rd_out_r1[247]
  PIN rd_out_r1[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 481.285 0.070 481.355 ;
    END
  END rd_out_r1[248]
  PIN rd_out_r1[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 481.845 0.070 481.915 ;
    END
  END rd_out_r1[249]
  PIN rd_out_r1[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 482.405 0.070 482.475 ;
    END
  END rd_out_r1[250]
  PIN rd_out_r1[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 482.965 0.070 483.035 ;
    END
  END rd_out_r1[251]
  PIN rd_out_r1[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 483.525 0.070 483.595 ;
    END
  END rd_out_r1[252]
  PIN rd_out_r1[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 484.085 0.070 484.155 ;
    END
  END rd_out_r1[253]
  PIN rd_out_r1[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 484.645 0.070 484.715 ;
    END
  END rd_out_r1[254]
  PIN rd_out_r1[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 485.205 0.070 485.275 ;
    END
  END rd_out_r1[255]
  PIN rd_out_r1[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 485.765 0.070 485.835 ;
    END
  END rd_out_r1[256]
  PIN rd_out_r1[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 486.325 0.070 486.395 ;
    END
  END rd_out_r1[257]
  PIN rd_out_r1[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 486.885 0.070 486.955 ;
    END
  END rd_out_r1[258]
  PIN rd_out_r1[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 487.445 0.070 487.515 ;
    END
  END rd_out_r1[259]
  PIN rd_out_r1[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 488.005 0.070 488.075 ;
    END
  END rd_out_r1[260]
  PIN rd_out_r1[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 488.565 0.070 488.635 ;
    END
  END rd_out_r1[261]
  PIN rd_out_r1[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 489.125 0.070 489.195 ;
    END
  END rd_out_r1[262]
  PIN rd_out_r1[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 489.685 0.070 489.755 ;
    END
  END rd_out_r1[263]
  PIN rd_out_r1[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 490.245 0.070 490.315 ;
    END
  END rd_out_r1[264]
  PIN rd_out_r1[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 490.805 0.070 490.875 ;
    END
  END rd_out_r1[265]
  PIN rd_out_r1[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 491.365 0.070 491.435 ;
    END
  END rd_out_r1[266]
  PIN rd_out_r1[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 491.925 0.070 491.995 ;
    END
  END rd_out_r1[267]
  PIN rd_out_r1[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 492.485 0.070 492.555 ;
    END
  END rd_out_r1[268]
  PIN rd_out_r1[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 493.045 0.070 493.115 ;
    END
  END rd_out_r1[269]
  PIN rd_out_r1[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 493.605 0.070 493.675 ;
    END
  END rd_out_r1[270]
  PIN rd_out_r1[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 494.165 0.070 494.235 ;
    END
  END rd_out_r1[271]
  PIN rd_out_r1[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 494.725 0.070 494.795 ;
    END
  END rd_out_r1[272]
  PIN rd_out_r1[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 495.285 0.070 495.355 ;
    END
  END rd_out_r1[273]
  PIN rd_out_r1[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 495.845 0.070 495.915 ;
    END
  END rd_out_r1[274]
  PIN rd_out_r1[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 496.405 0.070 496.475 ;
    END
  END rd_out_r1[275]
  PIN rd_out_r1[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 496.965 0.070 497.035 ;
    END
  END rd_out_r1[276]
  PIN rd_out_r1[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 497.525 0.070 497.595 ;
    END
  END rd_out_r1[277]
  PIN rd_out_r1[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 498.085 0.070 498.155 ;
    END
  END rd_out_r1[278]
  PIN rd_out_r1[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 498.645 0.070 498.715 ;
    END
  END rd_out_r1[279]
  PIN rd_out_r1[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 499.205 0.070 499.275 ;
    END
  END rd_out_r1[280]
  PIN rd_out_r1[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 499.765 0.070 499.835 ;
    END
  END rd_out_r1[281]
  PIN rd_out_r1[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 500.325 0.070 500.395 ;
    END
  END rd_out_r1[282]
  PIN rd_out_r1[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 500.885 0.070 500.955 ;
    END
  END rd_out_r1[283]
  PIN rd_out_r1[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 501.445 0.070 501.515 ;
    END
  END rd_out_r1[284]
  PIN rd_out_r1[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 502.005 0.070 502.075 ;
    END
  END rd_out_r1[285]
  PIN rd_out_r1[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 502.565 0.070 502.635 ;
    END
  END rd_out_r1[286]
  PIN rd_out_r1[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 503.125 0.070 503.195 ;
    END
  END rd_out_r1[287]
  PIN rd_out_r1[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 503.685 0.070 503.755 ;
    END
  END rd_out_r1[288]
  PIN rd_out_r1[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 504.245 0.070 504.315 ;
    END
  END rd_out_r1[289]
  PIN rd_out_r1[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 504.805 0.070 504.875 ;
    END
  END rd_out_r1[290]
  PIN rd_out_r1[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.365 0.070 505.435 ;
    END
  END rd_out_r1[291]
  PIN rd_out_r1[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.925 0.070 505.995 ;
    END
  END rd_out_r1[292]
  PIN rd_out_r1[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 506.485 0.070 506.555 ;
    END
  END rd_out_r1[293]
  PIN rd_out_r1[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.045 0.070 507.115 ;
    END
  END rd_out_r1[294]
  PIN rd_out_r1[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.605 0.070 507.675 ;
    END
  END rd_out_r1[295]
  PIN rd_out_r1[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 508.165 0.070 508.235 ;
    END
  END rd_out_r1[296]
  PIN rd_out_r1[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 508.725 0.070 508.795 ;
    END
  END rd_out_r1[297]
  PIN rd_out_r1[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.285 0.070 509.355 ;
    END
  END rd_out_r1[298]
  PIN rd_out_r1[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.845 0.070 509.915 ;
    END
  END rd_out_r1[299]
  PIN rd_out_r1[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.405 0.070 510.475 ;
    END
  END rd_out_r1[300]
  PIN rd_out_r1[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.965 0.070 511.035 ;
    END
  END rd_out_r1[301]
  PIN rd_out_r1[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 511.525 0.070 511.595 ;
    END
  END rd_out_r1[302]
  PIN rd_out_r1[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.085 0.070 512.155 ;
    END
  END rd_out_r1[303]
  PIN rd_out_r1[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.645 0.070 512.715 ;
    END
  END rd_out_r1[304]
  PIN rd_out_r1[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 513.205 0.070 513.275 ;
    END
  END rd_out_r1[305]
  PIN rd_out_r1[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 513.765 0.070 513.835 ;
    END
  END rd_out_r1[306]
  PIN rd_out_r1[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.325 0.070 514.395 ;
    END
  END rd_out_r1[307]
  PIN rd_out_r1[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.885 0.070 514.955 ;
    END
  END rd_out_r1[308]
  PIN rd_out_r1[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 515.445 0.070 515.515 ;
    END
  END rd_out_r1[309]
  PIN rd_out_r1[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.005 0.070 516.075 ;
    END
  END rd_out_r1[310]
  PIN rd_out_r1[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.565 0.070 516.635 ;
    END
  END rd_out_r1[311]
  PIN rd_out_r1[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.125 0.070 517.195 ;
    END
  END rd_out_r1[312]
  PIN rd_out_r1[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.685 0.070 517.755 ;
    END
  END rd_out_r1[313]
  PIN rd_out_r1[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.245 0.070 518.315 ;
    END
  END rd_out_r1[314]
  PIN rd_out_r1[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.805 0.070 518.875 ;
    END
  END rd_out_r1[315]
  PIN rd_out_r1[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.365 0.070 519.435 ;
    END
  END rd_out_r1[316]
  PIN rd_out_r1[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.925 0.070 519.995 ;
    END
  END rd_out_r1[317]
  PIN rd_out_r1[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.485 0.070 520.555 ;
    END
  END rd_out_r1[318]
  PIN rd_out_r1[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.045 0.070 521.115 ;
    END
  END rd_out_r1[319]
  PIN rd_out_r1[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.605 0.070 521.675 ;
    END
  END rd_out_r1[320]
  PIN rd_out_r1[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.165 0.070 522.235 ;
    END
  END rd_out_r1[321]
  PIN rd_out_r1[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.725 0.070 522.795 ;
    END
  END rd_out_r1[322]
  PIN rd_out_r1[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.285 0.070 523.355 ;
    END
  END rd_out_r1[323]
  PIN rd_out_r1[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.845 0.070 523.915 ;
    END
  END rd_out_r1[324]
  PIN rd_out_r1[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.405 0.070 524.475 ;
    END
  END rd_out_r1[325]
  PIN rd_out_r1[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.965 0.070 525.035 ;
    END
  END rd_out_r1[326]
  PIN rd_out_r1[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.525 0.070 525.595 ;
    END
  END rd_out_r1[327]
  PIN rd_out_r1[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.085 0.070 526.155 ;
    END
  END rd_out_r1[328]
  PIN rd_out_r1[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.645 0.070 526.715 ;
    END
  END rd_out_r1[329]
  PIN rd_out_r1[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.205 0.070 527.275 ;
    END
  END rd_out_r1[330]
  PIN rd_out_r1[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.765 0.070 527.835 ;
    END
  END rd_out_r1[331]
  PIN rd_out_r1[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.325 0.070 528.395 ;
    END
  END rd_out_r1[332]
  PIN rd_out_r1[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.885 0.070 528.955 ;
    END
  END rd_out_r1[333]
  PIN rd_out_r1[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.445 0.070 529.515 ;
    END
  END rd_out_r1[334]
  PIN rd_out_r1[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.005 0.070 530.075 ;
    END
  END rd_out_r1[335]
  PIN rd_out_r1[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.565 0.070 530.635 ;
    END
  END rd_out_r1[336]
  PIN rd_out_r1[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.125 0.070 531.195 ;
    END
  END rd_out_r1[337]
  PIN rd_out_r1[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.685 0.070 531.755 ;
    END
  END rd_out_r1[338]
  PIN rd_out_r1[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.245 0.070 532.315 ;
    END
  END rd_out_r1[339]
  PIN rd_out_r1[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.805 0.070 532.875 ;
    END
  END rd_out_r1[340]
  PIN rd_out_r1[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.365 0.070 533.435 ;
    END
  END rd_out_r1[341]
  PIN rd_out_r1[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.925 0.070 533.995 ;
    END
  END rd_out_r1[342]
  PIN rd_out_r1[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.485 0.070 534.555 ;
    END
  END rd_out_r1[343]
  PIN rd_out_r1[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.045 0.070 535.115 ;
    END
  END rd_out_r1[344]
  PIN rd_out_r1[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.605 0.070 535.675 ;
    END
  END rd_out_r1[345]
  PIN rd_out_r1[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.165 0.070 536.235 ;
    END
  END rd_out_r1[346]
  PIN rd_out_r1[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.725 0.070 536.795 ;
    END
  END rd_out_r1[347]
  PIN rd_out_r1[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.285 0.070 537.355 ;
    END
  END rd_out_r1[348]
  PIN rd_out_r1[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.845 0.070 537.915 ;
    END
  END rd_out_r1[349]
  PIN rd_out_r1[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.405 0.070 538.475 ;
    END
  END rd_out_r1[350]
  PIN rd_out_r1[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.965 0.070 539.035 ;
    END
  END rd_out_r1[351]
  PIN rd_out_r1[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.525 0.070 539.595 ;
    END
  END rd_out_r1[352]
  PIN rd_out_r1[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.085 0.070 540.155 ;
    END
  END rd_out_r1[353]
  PIN rd_out_r1[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.645 0.070 540.715 ;
    END
  END rd_out_r1[354]
  PIN rd_out_r1[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.205 0.070 541.275 ;
    END
  END rd_out_r1[355]
  PIN rd_out_r1[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.765 0.070 541.835 ;
    END
  END rd_out_r1[356]
  PIN rd_out_r1[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.325 0.070 542.395 ;
    END
  END rd_out_r1[357]
  PIN rd_out_r1[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.885 0.070 542.955 ;
    END
  END rd_out_r1[358]
  PIN rd_out_r1[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.445 0.070 543.515 ;
    END
  END rd_out_r1[359]
  PIN rd_out_r1[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.005 0.070 544.075 ;
    END
  END rd_out_r1[360]
  PIN rd_out_r1[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.565 0.070 544.635 ;
    END
  END rd_out_r1[361]
  PIN rd_out_r1[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.125 0.070 545.195 ;
    END
  END rd_out_r1[362]
  PIN rd_out_r1[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.685 0.070 545.755 ;
    END
  END rd_out_r1[363]
  PIN rd_out_r1[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.245 0.070 546.315 ;
    END
  END rd_out_r1[364]
  PIN rd_out_r1[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.805 0.070 546.875 ;
    END
  END rd_out_r1[365]
  PIN rd_out_r1[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.365 0.070 547.435 ;
    END
  END rd_out_r1[366]
  PIN rd_out_r1[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.925 0.070 547.995 ;
    END
  END rd_out_r1[367]
  PIN rd_out_r1[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.485 0.070 548.555 ;
    END
  END rd_out_r1[368]
  PIN rd_out_r1[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.045 0.070 549.115 ;
    END
  END rd_out_r1[369]
  PIN rd_out_r1[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.605 0.070 549.675 ;
    END
  END rd_out_r1[370]
  PIN rd_out_r1[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.165 0.070 550.235 ;
    END
  END rd_out_r1[371]
  PIN rd_out_r1[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.725 0.070 550.795 ;
    END
  END rd_out_r1[372]
  PIN rd_out_r1[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.285 0.070 551.355 ;
    END
  END rd_out_r1[373]
  PIN rd_out_r1[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.845 0.070 551.915 ;
    END
  END rd_out_r1[374]
  PIN rd_out_r1[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.405 0.070 552.475 ;
    END
  END rd_out_r1[375]
  PIN rd_out_r1[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.965 0.070 553.035 ;
    END
  END rd_out_r1[376]
  PIN rd_out_r1[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.525 0.070 553.595 ;
    END
  END rd_out_r1[377]
  PIN rd_out_r1[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.085 0.070 554.155 ;
    END
  END rd_out_r1[378]
  PIN rd_out_r1[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.645 0.070 554.715 ;
    END
  END rd_out_r1[379]
  PIN rd_out_r1[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.205 0.070 555.275 ;
    END
  END rd_out_r1[380]
  PIN rd_out_r1[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.765 0.070 555.835 ;
    END
  END rd_out_r1[381]
  PIN rd_out_r1[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.325 0.070 556.395 ;
    END
  END rd_out_r1[382]
  PIN rd_out_r1[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.885 0.070 556.955 ;
    END
  END rd_out_r1[383]
  PIN rd_out_r1[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.445 0.070 557.515 ;
    END
  END rd_out_r1[384]
  PIN rd_out_r1[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.005 0.070 558.075 ;
    END
  END rd_out_r1[385]
  PIN rd_out_r1[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.565 0.070 558.635 ;
    END
  END rd_out_r1[386]
  PIN rd_out_r1[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.125 0.070 559.195 ;
    END
  END rd_out_r1[387]
  PIN rd_out_r1[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.685 0.070 559.755 ;
    END
  END rd_out_r1[388]
  PIN rd_out_r1[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.245 0.070 560.315 ;
    END
  END rd_out_r1[389]
  PIN rd_out_r1[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.805 0.070 560.875 ;
    END
  END rd_out_r1[390]
  PIN rd_out_r1[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.365 0.070 561.435 ;
    END
  END rd_out_r1[391]
  PIN rd_out_r1[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.925 0.070 561.995 ;
    END
  END rd_out_r1[392]
  PIN rd_out_r1[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.485 0.070 562.555 ;
    END
  END rd_out_r1[393]
  PIN rd_out_r1[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.045 0.070 563.115 ;
    END
  END rd_out_r1[394]
  PIN rd_out_r1[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.605 0.070 563.675 ;
    END
  END rd_out_r1[395]
  PIN rd_out_r1[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.165 0.070 564.235 ;
    END
  END rd_out_r1[396]
  PIN rd_out_r1[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.725 0.070 564.795 ;
    END
  END rd_out_r1[397]
  PIN rd_out_r1[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.285 0.070 565.355 ;
    END
  END rd_out_r1[398]
  PIN rd_out_r1[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.845 0.070 565.915 ;
    END
  END rd_out_r1[399]
  PIN rd_out_r1[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.405 0.070 566.475 ;
    END
  END rd_out_r1[400]
  PIN rd_out_r1[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.965 0.070 567.035 ;
    END
  END rd_out_r1[401]
  PIN rd_out_r1[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.525 0.070 567.595 ;
    END
  END rd_out_r1[402]
  PIN rd_out_r1[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.085 0.070 568.155 ;
    END
  END rd_out_r1[403]
  PIN rd_out_r1[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.645 0.070 568.715 ;
    END
  END rd_out_r1[404]
  PIN rd_out_r1[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.205 0.070 569.275 ;
    END
  END rd_out_r1[405]
  PIN rd_out_r1[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.765 0.070 569.835 ;
    END
  END rd_out_r1[406]
  PIN rd_out_r1[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.325 0.070 570.395 ;
    END
  END rd_out_r1[407]
  PIN rd_out_r1[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.885 0.070 570.955 ;
    END
  END rd_out_r1[408]
  PIN rd_out_r1[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.445 0.070 571.515 ;
    END
  END rd_out_r1[409]
  PIN rd_out_r1[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.005 0.070 572.075 ;
    END
  END rd_out_r1[410]
  PIN rd_out_r1[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.565 0.070 572.635 ;
    END
  END rd_out_r1[411]
  PIN rd_out_r1[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.125 0.070 573.195 ;
    END
  END rd_out_r1[412]
  PIN rd_out_r1[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.685 0.070 573.755 ;
    END
  END rd_out_r1[413]
  PIN rd_out_r1[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.245 0.070 574.315 ;
    END
  END rd_out_r1[414]
  PIN rd_out_r1[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.805 0.070 574.875 ;
    END
  END rd_out_r1[415]
  PIN rd_out_r1[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.365 0.070 575.435 ;
    END
  END rd_out_r1[416]
  PIN rd_out_r1[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.925 0.070 575.995 ;
    END
  END rd_out_r1[417]
  PIN rd_out_r1[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 576.485 0.070 576.555 ;
    END
  END rd_out_r1[418]
  PIN rd_out_r1[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.045 0.070 577.115 ;
    END
  END rd_out_r1[419]
  PIN rd_out_r1[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.605 0.070 577.675 ;
    END
  END rd_out_r1[420]
  PIN rd_out_r1[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.165 0.070 578.235 ;
    END
  END rd_out_r1[421]
  PIN rd_out_r1[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.725 0.070 578.795 ;
    END
  END rd_out_r1[422]
  PIN rd_out_r1[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.285 0.070 579.355 ;
    END
  END rd_out_r1[423]
  PIN rd_out_r1[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.845 0.070 579.915 ;
    END
  END rd_out_r1[424]
  PIN rd_out_r1[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.405 0.070 580.475 ;
    END
  END rd_out_r1[425]
  PIN rd_out_r1[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.965 0.070 581.035 ;
    END
  END rd_out_r1[426]
  PIN rd_out_r1[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 581.525 0.070 581.595 ;
    END
  END rd_out_r1[427]
  PIN rd_out_r1[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.085 0.070 582.155 ;
    END
  END rd_out_r1[428]
  PIN rd_out_r1[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.645 0.070 582.715 ;
    END
  END rd_out_r1[429]
  PIN rd_out_r1[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.205 0.070 583.275 ;
    END
  END rd_out_r1[430]
  PIN rd_out_r1[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.765 0.070 583.835 ;
    END
  END rd_out_r1[431]
  PIN rd_out_r1[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.325 0.070 584.395 ;
    END
  END rd_out_r1[432]
  PIN rd_out_r1[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.885 0.070 584.955 ;
    END
  END rd_out_r1[433]
  PIN rd_out_r1[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 585.445 0.070 585.515 ;
    END
  END rd_out_r1[434]
  PIN rd_out_r1[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.005 0.070 586.075 ;
    END
  END rd_out_r1[435]
  PIN rd_out_r1[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.565 0.070 586.635 ;
    END
  END rd_out_r1[436]
  PIN rd_out_r1[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.125 0.070 587.195 ;
    END
  END rd_out_r1[437]
  PIN rd_out_r1[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.685 0.070 587.755 ;
    END
  END rd_out_r1[438]
  PIN rd_out_r1[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.245 0.070 588.315 ;
    END
  END rd_out_r1[439]
  PIN rd_out_r1[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.805 0.070 588.875 ;
    END
  END rd_out_r1[440]
  PIN rd_out_r1[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.365 0.070 589.435 ;
    END
  END rd_out_r1[441]
  PIN rd_out_r1[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.925 0.070 589.995 ;
    END
  END rd_out_r1[442]
  PIN rd_out_r1[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 590.485 0.070 590.555 ;
    END
  END rd_out_r1[443]
  PIN rd_out_r1[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.045 0.070 591.115 ;
    END
  END rd_out_r1[444]
  PIN rd_out_r1[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.605 0.070 591.675 ;
    END
  END rd_out_r1[445]
  PIN rd_out_r1[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.165 0.070 592.235 ;
    END
  END rd_out_r1[446]
  PIN rd_out_r1[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.725 0.070 592.795 ;
    END
  END rd_out_r1[447]
  PIN rd_out_r1[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.285 0.070 593.355 ;
    END
  END rd_out_r1[448]
  PIN rd_out_r1[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.845 0.070 593.915 ;
    END
  END rd_out_r1[449]
  PIN rd_out_r1[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.405 0.070 594.475 ;
    END
  END rd_out_r1[450]
  PIN rd_out_r1[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.965 0.070 595.035 ;
    END
  END rd_out_r1[451]
  PIN rd_out_r1[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.525 0.070 595.595 ;
    END
  END rd_out_r1[452]
  PIN rd_out_r1[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.085 0.070 596.155 ;
    END
  END rd_out_r1[453]
  PIN rd_out_r1[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.645 0.070 596.715 ;
    END
  END rd_out_r1[454]
  PIN rd_out_r1[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.205 0.070 597.275 ;
    END
  END rd_out_r1[455]
  PIN rd_out_r1[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.765 0.070 597.835 ;
    END
  END rd_out_r1[456]
  PIN rd_out_r1[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.325 0.070 598.395 ;
    END
  END rd_out_r1[457]
  PIN rd_out_r1[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.885 0.070 598.955 ;
    END
  END rd_out_r1[458]
  PIN rd_out_r1[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.445 0.070 599.515 ;
    END
  END rd_out_r1[459]
  PIN rd_out_r1[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.005 0.070 600.075 ;
    END
  END rd_out_r1[460]
  PIN rd_out_r1[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.565 0.070 600.635 ;
    END
  END rd_out_r1[461]
  PIN rd_out_r1[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.125 0.070 601.195 ;
    END
  END rd_out_r1[462]
  PIN rd_out_r1[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.685 0.070 601.755 ;
    END
  END rd_out_r1[463]
  PIN rd_out_r1[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.245 0.070 602.315 ;
    END
  END rd_out_r1[464]
  PIN rd_out_r1[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.805 0.070 602.875 ;
    END
  END rd_out_r1[465]
  PIN rd_out_r1[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.365 0.070 603.435 ;
    END
  END rd_out_r1[466]
  PIN rd_out_r1[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.925 0.070 603.995 ;
    END
  END rd_out_r1[467]
  PIN rd_out_r1[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.485 0.070 604.555 ;
    END
  END rd_out_r1[468]
  PIN rd_out_r1[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.045 0.070 605.115 ;
    END
  END rd_out_r1[469]
  PIN rd_out_r1[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.605 0.070 605.675 ;
    END
  END rd_out_r1[470]
  PIN rd_out_r1[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.165 0.070 606.235 ;
    END
  END rd_out_r1[471]
  PIN rd_out_r1[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.725 0.070 606.795 ;
    END
  END rd_out_r1[472]
  PIN rd_out_r1[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.285 0.070 607.355 ;
    END
  END rd_out_r1[473]
  PIN rd_out_r1[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.845 0.070 607.915 ;
    END
  END rd_out_r1[474]
  PIN rd_out_r1[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.405 0.070 608.475 ;
    END
  END rd_out_r1[475]
  PIN rd_out_r1[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.965 0.070 609.035 ;
    END
  END rd_out_r1[476]
  PIN rd_out_r1[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.525 0.070 609.595 ;
    END
  END rd_out_r1[477]
  PIN rd_out_r1[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.085 0.070 610.155 ;
    END
  END rd_out_r1[478]
  PIN rd_out_r1[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.645 0.070 610.715 ;
    END
  END rd_out_r1[479]
  PIN rd_out_r1[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.205 0.070 611.275 ;
    END
  END rd_out_r1[480]
  PIN rd_out_r1[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.765 0.070 611.835 ;
    END
  END rd_out_r1[481]
  PIN rd_out_r1[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.325 0.070 612.395 ;
    END
  END rd_out_r1[482]
  PIN rd_out_r1[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.885 0.070 612.955 ;
    END
  END rd_out_r1[483]
  PIN rd_out_r1[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 613.445 0.070 613.515 ;
    END
  END rd_out_r1[484]
  PIN rd_out_r1[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.005 0.070 614.075 ;
    END
  END rd_out_r1[485]
  PIN rd_out_r1[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.565 0.070 614.635 ;
    END
  END rd_out_r1[486]
  PIN rd_out_r1[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.125 0.070 615.195 ;
    END
  END rd_out_r1[487]
  PIN rd_out_r1[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.685 0.070 615.755 ;
    END
  END rd_out_r1[488]
  PIN rd_out_r1[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.245 0.070 616.315 ;
    END
  END rd_out_r1[489]
  PIN rd_out_r1[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.805 0.070 616.875 ;
    END
  END rd_out_r1[490]
  PIN rd_out_r1[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.365 0.070 617.435 ;
    END
  END rd_out_r1[491]
  PIN rd_out_r1[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.925 0.070 617.995 ;
    END
  END rd_out_r1[492]
  PIN rd_out_r1[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.485 0.070 618.555 ;
    END
  END rd_out_r1[493]
  PIN rd_out_r1[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.045 0.070 619.115 ;
    END
  END rd_out_r1[494]
  PIN rd_out_r1[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.605 0.070 619.675 ;
    END
  END rd_out_r1[495]
  PIN rd_out_r1[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.165 0.070 620.235 ;
    END
  END rd_out_r1[496]
  PIN rd_out_r1[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.725 0.070 620.795 ;
    END
  END rd_out_r1[497]
  PIN rd_out_r1[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.285 0.070 621.355 ;
    END
  END rd_out_r1[498]
  PIN rd_out_r1[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.845 0.070 621.915 ;
    END
  END rd_out_r1[499]
  PIN rd_out_r1[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.405 0.070 622.475 ;
    END
  END rd_out_r1[500]
  PIN rd_out_r1[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.965 0.070 623.035 ;
    END
  END rd_out_r1[501]
  PIN rd_out_r1[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.525 0.070 623.595 ;
    END
  END rd_out_r1[502]
  PIN rd_out_r1[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.085 0.070 624.155 ;
    END
  END rd_out_r1[503]
  PIN rd_out_r1[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.645 0.070 624.715 ;
    END
  END rd_out_r1[504]
  PIN rd_out_r1[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.205 0.070 625.275 ;
    END
  END rd_out_r1[505]
  PIN rd_out_r1[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.765 0.070 625.835 ;
    END
  END rd_out_r1[506]
  PIN rd_out_r1[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.325 0.070 626.395 ;
    END
  END rd_out_r1[507]
  PIN rd_out_r1[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.885 0.070 626.955 ;
    END
  END rd_out_r1[508]
  PIN rd_out_r1[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 627.445 0.070 627.515 ;
    END
  END rd_out_r1[509]
  PIN rd_out_r1[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.005 0.070 628.075 ;
    END
  END rd_out_r1[510]
  PIN rd_out_r1[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.565 0.070 628.635 ;
    END
  END rd_out_r1[511]
  PIN wd_in_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.285 0.070 656.355 ;
    END
  END wd_in_w1[0]
  PIN wd_in_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.845 0.070 656.915 ;
    END
  END wd_in_w1[1]
  PIN wd_in_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.405 0.070 657.475 ;
    END
  END wd_in_w1[2]
  PIN wd_in_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.965 0.070 658.035 ;
    END
  END wd_in_w1[3]
  PIN wd_in_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.525 0.070 658.595 ;
    END
  END wd_in_w1[4]
  PIN wd_in_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.085 0.070 659.155 ;
    END
  END wd_in_w1[5]
  PIN wd_in_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.645 0.070 659.715 ;
    END
  END wd_in_w1[6]
  PIN wd_in_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.205 0.070 660.275 ;
    END
  END wd_in_w1[7]
  PIN wd_in_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.765 0.070 660.835 ;
    END
  END wd_in_w1[8]
  PIN wd_in_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.325 0.070 661.395 ;
    END
  END wd_in_w1[9]
  PIN wd_in_w1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.885 0.070 661.955 ;
    END
  END wd_in_w1[10]
  PIN wd_in_w1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.445 0.070 662.515 ;
    END
  END wd_in_w1[11]
  PIN wd_in_w1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.005 0.070 663.075 ;
    END
  END wd_in_w1[12]
  PIN wd_in_w1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.565 0.070 663.635 ;
    END
  END wd_in_w1[13]
  PIN wd_in_w1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.125 0.070 664.195 ;
    END
  END wd_in_w1[14]
  PIN wd_in_w1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.685 0.070 664.755 ;
    END
  END wd_in_w1[15]
  PIN wd_in_w1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.245 0.070 665.315 ;
    END
  END wd_in_w1[16]
  PIN wd_in_w1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.805 0.070 665.875 ;
    END
  END wd_in_w1[17]
  PIN wd_in_w1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.365 0.070 666.435 ;
    END
  END wd_in_w1[18]
  PIN wd_in_w1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.925 0.070 666.995 ;
    END
  END wd_in_w1[19]
  PIN wd_in_w1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.485 0.070 667.555 ;
    END
  END wd_in_w1[20]
  PIN wd_in_w1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.045 0.070 668.115 ;
    END
  END wd_in_w1[21]
  PIN wd_in_w1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.605 0.070 668.675 ;
    END
  END wd_in_w1[22]
  PIN wd_in_w1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.165 0.070 669.235 ;
    END
  END wd_in_w1[23]
  PIN wd_in_w1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.725 0.070 669.795 ;
    END
  END wd_in_w1[24]
  PIN wd_in_w1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.285 0.070 670.355 ;
    END
  END wd_in_w1[25]
  PIN wd_in_w1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.845 0.070 670.915 ;
    END
  END wd_in_w1[26]
  PIN wd_in_w1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.405 0.070 671.475 ;
    END
  END wd_in_w1[27]
  PIN wd_in_w1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.965 0.070 672.035 ;
    END
  END wd_in_w1[28]
  PIN wd_in_w1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.525 0.070 672.595 ;
    END
  END wd_in_w1[29]
  PIN wd_in_w1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.085 0.070 673.155 ;
    END
  END wd_in_w1[30]
  PIN wd_in_w1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.645 0.070 673.715 ;
    END
  END wd_in_w1[31]
  PIN wd_in_w1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.205 0.070 674.275 ;
    END
  END wd_in_w1[32]
  PIN wd_in_w1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.765 0.070 674.835 ;
    END
  END wd_in_w1[33]
  PIN wd_in_w1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.325 0.070 675.395 ;
    END
  END wd_in_w1[34]
  PIN wd_in_w1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.885 0.070 675.955 ;
    END
  END wd_in_w1[35]
  PIN wd_in_w1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 676.445 0.070 676.515 ;
    END
  END wd_in_w1[36]
  PIN wd_in_w1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.005 0.070 677.075 ;
    END
  END wd_in_w1[37]
  PIN wd_in_w1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.565 0.070 677.635 ;
    END
  END wd_in_w1[38]
  PIN wd_in_w1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.125 0.070 678.195 ;
    END
  END wd_in_w1[39]
  PIN wd_in_w1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.685 0.070 678.755 ;
    END
  END wd_in_w1[40]
  PIN wd_in_w1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.245 0.070 679.315 ;
    END
  END wd_in_w1[41]
  PIN wd_in_w1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.805 0.070 679.875 ;
    END
  END wd_in_w1[42]
  PIN wd_in_w1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.365 0.070 680.435 ;
    END
  END wd_in_w1[43]
  PIN wd_in_w1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.925 0.070 680.995 ;
    END
  END wd_in_w1[44]
  PIN wd_in_w1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.485 0.070 681.555 ;
    END
  END wd_in_w1[45]
  PIN wd_in_w1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.045 0.070 682.115 ;
    END
  END wd_in_w1[46]
  PIN wd_in_w1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.605 0.070 682.675 ;
    END
  END wd_in_w1[47]
  PIN wd_in_w1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.165 0.070 683.235 ;
    END
  END wd_in_w1[48]
  PIN wd_in_w1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.725 0.070 683.795 ;
    END
  END wd_in_w1[49]
  PIN wd_in_w1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.285 0.070 684.355 ;
    END
  END wd_in_w1[50]
  PIN wd_in_w1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.845 0.070 684.915 ;
    END
  END wd_in_w1[51]
  PIN wd_in_w1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.405 0.070 685.475 ;
    END
  END wd_in_w1[52]
  PIN wd_in_w1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.965 0.070 686.035 ;
    END
  END wd_in_w1[53]
  PIN wd_in_w1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 686.525 0.070 686.595 ;
    END
  END wd_in_w1[54]
  PIN wd_in_w1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.085 0.070 687.155 ;
    END
  END wd_in_w1[55]
  PIN wd_in_w1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.645 0.070 687.715 ;
    END
  END wd_in_w1[56]
  PIN wd_in_w1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.205 0.070 688.275 ;
    END
  END wd_in_w1[57]
  PIN wd_in_w1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.765 0.070 688.835 ;
    END
  END wd_in_w1[58]
  PIN wd_in_w1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.325 0.070 689.395 ;
    END
  END wd_in_w1[59]
  PIN wd_in_w1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.885 0.070 689.955 ;
    END
  END wd_in_w1[60]
  PIN wd_in_w1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 690.445 0.070 690.515 ;
    END
  END wd_in_w1[61]
  PIN wd_in_w1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.005 0.070 691.075 ;
    END
  END wd_in_w1[62]
  PIN wd_in_w1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.565 0.070 691.635 ;
    END
  END wd_in_w1[63]
  PIN wd_in_w1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.125 0.070 692.195 ;
    END
  END wd_in_w1[64]
  PIN wd_in_w1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.685 0.070 692.755 ;
    END
  END wd_in_w1[65]
  PIN wd_in_w1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.245 0.070 693.315 ;
    END
  END wd_in_w1[66]
  PIN wd_in_w1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.805 0.070 693.875 ;
    END
  END wd_in_w1[67]
  PIN wd_in_w1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.365 0.070 694.435 ;
    END
  END wd_in_w1[68]
  PIN wd_in_w1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.925 0.070 694.995 ;
    END
  END wd_in_w1[69]
  PIN wd_in_w1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 695.485 0.070 695.555 ;
    END
  END wd_in_w1[70]
  PIN wd_in_w1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.045 0.070 696.115 ;
    END
  END wd_in_w1[71]
  PIN wd_in_w1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.605 0.070 696.675 ;
    END
  END wd_in_w1[72]
  PIN wd_in_w1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 697.165 0.070 697.235 ;
    END
  END wd_in_w1[73]
  PIN wd_in_w1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 697.725 0.070 697.795 ;
    END
  END wd_in_w1[74]
  PIN wd_in_w1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.285 0.070 698.355 ;
    END
  END wd_in_w1[75]
  PIN wd_in_w1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.845 0.070 698.915 ;
    END
  END wd_in_w1[76]
  PIN wd_in_w1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 699.405 0.070 699.475 ;
    END
  END wd_in_w1[77]
  PIN wd_in_w1[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 699.965 0.070 700.035 ;
    END
  END wd_in_w1[78]
  PIN wd_in_w1[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 700.525 0.070 700.595 ;
    END
  END wd_in_w1[79]
  PIN wd_in_w1[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.085 0.070 701.155 ;
    END
  END wd_in_w1[80]
  PIN wd_in_w1[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.645 0.070 701.715 ;
    END
  END wd_in_w1[81]
  PIN wd_in_w1[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.205 0.070 702.275 ;
    END
  END wd_in_w1[82]
  PIN wd_in_w1[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.765 0.070 702.835 ;
    END
  END wd_in_w1[83]
  PIN wd_in_w1[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.325 0.070 703.395 ;
    END
  END wd_in_w1[84]
  PIN wd_in_w1[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.885 0.070 703.955 ;
    END
  END wd_in_w1[85]
  PIN wd_in_w1[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.445 0.070 704.515 ;
    END
  END wd_in_w1[86]
  PIN wd_in_w1[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.005 0.070 705.075 ;
    END
  END wd_in_w1[87]
  PIN wd_in_w1[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.565 0.070 705.635 ;
    END
  END wd_in_w1[88]
  PIN wd_in_w1[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.125 0.070 706.195 ;
    END
  END wd_in_w1[89]
  PIN wd_in_w1[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.685 0.070 706.755 ;
    END
  END wd_in_w1[90]
  PIN wd_in_w1[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.245 0.070 707.315 ;
    END
  END wd_in_w1[91]
  PIN wd_in_w1[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.805 0.070 707.875 ;
    END
  END wd_in_w1[92]
  PIN wd_in_w1[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.365 0.070 708.435 ;
    END
  END wd_in_w1[93]
  PIN wd_in_w1[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.925 0.070 708.995 ;
    END
  END wd_in_w1[94]
  PIN wd_in_w1[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.485 0.070 709.555 ;
    END
  END wd_in_w1[95]
  PIN wd_in_w1[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.045 0.070 710.115 ;
    END
  END wd_in_w1[96]
  PIN wd_in_w1[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.605 0.070 710.675 ;
    END
  END wd_in_w1[97]
  PIN wd_in_w1[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 711.165 0.070 711.235 ;
    END
  END wd_in_w1[98]
  PIN wd_in_w1[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 711.725 0.070 711.795 ;
    END
  END wd_in_w1[99]
  PIN wd_in_w1[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.285 0.070 712.355 ;
    END
  END wd_in_w1[100]
  PIN wd_in_w1[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.845 0.070 712.915 ;
    END
  END wd_in_w1[101]
  PIN wd_in_w1[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 713.405 0.070 713.475 ;
    END
  END wd_in_w1[102]
  PIN wd_in_w1[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 713.965 0.070 714.035 ;
    END
  END wd_in_w1[103]
  PIN wd_in_w1[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 714.525 0.070 714.595 ;
    END
  END wd_in_w1[104]
  PIN wd_in_w1[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.085 0.070 715.155 ;
    END
  END wd_in_w1[105]
  PIN wd_in_w1[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.645 0.070 715.715 ;
    END
  END wd_in_w1[106]
  PIN wd_in_w1[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 716.205 0.070 716.275 ;
    END
  END wd_in_w1[107]
  PIN wd_in_w1[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 716.765 0.070 716.835 ;
    END
  END wd_in_w1[108]
  PIN wd_in_w1[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.325 0.070 717.395 ;
    END
  END wd_in_w1[109]
  PIN wd_in_w1[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.885 0.070 717.955 ;
    END
  END wd_in_w1[110]
  PIN wd_in_w1[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 718.445 0.070 718.515 ;
    END
  END wd_in_w1[111]
  PIN wd_in_w1[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.005 0.070 719.075 ;
    END
  END wd_in_w1[112]
  PIN wd_in_w1[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.565 0.070 719.635 ;
    END
  END wd_in_w1[113]
  PIN wd_in_w1[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 720.125 0.070 720.195 ;
    END
  END wd_in_w1[114]
  PIN wd_in_w1[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 720.685 0.070 720.755 ;
    END
  END wd_in_w1[115]
  PIN wd_in_w1[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.245 0.070 721.315 ;
    END
  END wd_in_w1[116]
  PIN wd_in_w1[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.805 0.070 721.875 ;
    END
  END wd_in_w1[117]
  PIN wd_in_w1[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.365 0.070 722.435 ;
    END
  END wd_in_w1[118]
  PIN wd_in_w1[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.925 0.070 722.995 ;
    END
  END wd_in_w1[119]
  PIN wd_in_w1[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.485 0.070 723.555 ;
    END
  END wd_in_w1[120]
  PIN wd_in_w1[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.045 0.070 724.115 ;
    END
  END wd_in_w1[121]
  PIN wd_in_w1[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.605 0.070 724.675 ;
    END
  END wd_in_w1[122]
  PIN wd_in_w1[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.165 0.070 725.235 ;
    END
  END wd_in_w1[123]
  PIN wd_in_w1[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.725 0.070 725.795 ;
    END
  END wd_in_w1[124]
  PIN wd_in_w1[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.285 0.070 726.355 ;
    END
  END wd_in_w1[125]
  PIN wd_in_w1[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.845 0.070 726.915 ;
    END
  END wd_in_w1[126]
  PIN wd_in_w1[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.405 0.070 727.475 ;
    END
  END wd_in_w1[127]
  PIN wd_in_w1[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.965 0.070 728.035 ;
    END
  END wd_in_w1[128]
  PIN wd_in_w1[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 728.525 0.070 728.595 ;
    END
  END wd_in_w1[129]
  PIN wd_in_w1[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.085 0.070 729.155 ;
    END
  END wd_in_w1[130]
  PIN wd_in_w1[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.645 0.070 729.715 ;
    END
  END wd_in_w1[131]
  PIN wd_in_w1[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.205 0.070 730.275 ;
    END
  END wd_in_w1[132]
  PIN wd_in_w1[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.765 0.070 730.835 ;
    END
  END wd_in_w1[133]
  PIN wd_in_w1[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 731.325 0.070 731.395 ;
    END
  END wd_in_w1[134]
  PIN wd_in_w1[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 731.885 0.070 731.955 ;
    END
  END wd_in_w1[135]
  PIN wd_in_w1[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 732.445 0.070 732.515 ;
    END
  END wd_in_w1[136]
  PIN wd_in_w1[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.005 0.070 733.075 ;
    END
  END wd_in_w1[137]
  PIN wd_in_w1[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.565 0.070 733.635 ;
    END
  END wd_in_w1[138]
  PIN wd_in_w1[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 734.125 0.070 734.195 ;
    END
  END wd_in_w1[139]
  PIN wd_in_w1[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 734.685 0.070 734.755 ;
    END
  END wd_in_w1[140]
  PIN wd_in_w1[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 735.245 0.070 735.315 ;
    END
  END wd_in_w1[141]
  PIN wd_in_w1[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 735.805 0.070 735.875 ;
    END
  END wd_in_w1[142]
  PIN wd_in_w1[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 736.365 0.070 736.435 ;
    END
  END wd_in_w1[143]
  PIN wd_in_w1[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 736.925 0.070 736.995 ;
    END
  END wd_in_w1[144]
  PIN wd_in_w1[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 737.485 0.070 737.555 ;
    END
  END wd_in_w1[145]
  PIN wd_in_w1[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 738.045 0.070 738.115 ;
    END
  END wd_in_w1[146]
  PIN wd_in_w1[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 738.605 0.070 738.675 ;
    END
  END wd_in_w1[147]
  PIN wd_in_w1[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 739.165 0.070 739.235 ;
    END
  END wd_in_w1[148]
  PIN wd_in_w1[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 739.725 0.070 739.795 ;
    END
  END wd_in_w1[149]
  PIN wd_in_w1[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.285 0.070 740.355 ;
    END
  END wd_in_w1[150]
  PIN wd_in_w1[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.845 0.070 740.915 ;
    END
  END wd_in_w1[151]
  PIN wd_in_w1[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 741.405 0.070 741.475 ;
    END
  END wd_in_w1[152]
  PIN wd_in_w1[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 741.965 0.070 742.035 ;
    END
  END wd_in_w1[153]
  PIN wd_in_w1[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 742.525 0.070 742.595 ;
    END
  END wd_in_w1[154]
  PIN wd_in_w1[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 743.085 0.070 743.155 ;
    END
  END wd_in_w1[155]
  PIN wd_in_w1[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 743.645 0.070 743.715 ;
    END
  END wd_in_w1[156]
  PIN wd_in_w1[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 744.205 0.070 744.275 ;
    END
  END wd_in_w1[157]
  PIN wd_in_w1[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 744.765 0.070 744.835 ;
    END
  END wd_in_w1[158]
  PIN wd_in_w1[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 745.325 0.070 745.395 ;
    END
  END wd_in_w1[159]
  PIN wd_in_w1[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 745.885 0.070 745.955 ;
    END
  END wd_in_w1[160]
  PIN wd_in_w1[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 746.445 0.070 746.515 ;
    END
  END wd_in_w1[161]
  PIN wd_in_w1[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.005 0.070 747.075 ;
    END
  END wd_in_w1[162]
  PIN wd_in_w1[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.565 0.070 747.635 ;
    END
  END wd_in_w1[163]
  PIN wd_in_w1[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 748.125 0.070 748.195 ;
    END
  END wd_in_w1[164]
  PIN wd_in_w1[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 748.685 0.070 748.755 ;
    END
  END wd_in_w1[165]
  PIN wd_in_w1[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 749.245 0.070 749.315 ;
    END
  END wd_in_w1[166]
  PIN wd_in_w1[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 749.805 0.070 749.875 ;
    END
  END wd_in_w1[167]
  PIN wd_in_w1[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 750.365 0.070 750.435 ;
    END
  END wd_in_w1[168]
  PIN wd_in_w1[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 750.925 0.070 750.995 ;
    END
  END wd_in_w1[169]
  PIN wd_in_w1[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 751.485 0.070 751.555 ;
    END
  END wd_in_w1[170]
  PIN wd_in_w1[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 752.045 0.070 752.115 ;
    END
  END wd_in_w1[171]
  PIN wd_in_w1[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 752.605 0.070 752.675 ;
    END
  END wd_in_w1[172]
  PIN wd_in_w1[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 753.165 0.070 753.235 ;
    END
  END wd_in_w1[173]
  PIN wd_in_w1[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 753.725 0.070 753.795 ;
    END
  END wd_in_w1[174]
  PIN wd_in_w1[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 754.285 0.070 754.355 ;
    END
  END wd_in_w1[175]
  PIN wd_in_w1[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 754.845 0.070 754.915 ;
    END
  END wd_in_w1[176]
  PIN wd_in_w1[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 755.405 0.070 755.475 ;
    END
  END wd_in_w1[177]
  PIN wd_in_w1[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 755.965 0.070 756.035 ;
    END
  END wd_in_w1[178]
  PIN wd_in_w1[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 756.525 0.070 756.595 ;
    END
  END wd_in_w1[179]
  PIN wd_in_w1[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 757.085 0.070 757.155 ;
    END
  END wd_in_w1[180]
  PIN wd_in_w1[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 757.645 0.070 757.715 ;
    END
  END wd_in_w1[181]
  PIN wd_in_w1[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 758.205 0.070 758.275 ;
    END
  END wd_in_w1[182]
  PIN wd_in_w1[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 758.765 0.070 758.835 ;
    END
  END wd_in_w1[183]
  PIN wd_in_w1[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.325 0.070 759.395 ;
    END
  END wd_in_w1[184]
  PIN wd_in_w1[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.885 0.070 759.955 ;
    END
  END wd_in_w1[185]
  PIN wd_in_w1[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 760.445 0.070 760.515 ;
    END
  END wd_in_w1[186]
  PIN wd_in_w1[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.005 0.070 761.075 ;
    END
  END wd_in_w1[187]
  PIN wd_in_w1[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.565 0.070 761.635 ;
    END
  END wd_in_w1[188]
  PIN wd_in_w1[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 762.125 0.070 762.195 ;
    END
  END wd_in_w1[189]
  PIN wd_in_w1[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 762.685 0.070 762.755 ;
    END
  END wd_in_w1[190]
  PIN wd_in_w1[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 763.245 0.070 763.315 ;
    END
  END wd_in_w1[191]
  PIN wd_in_w1[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 763.805 0.070 763.875 ;
    END
  END wd_in_w1[192]
  PIN wd_in_w1[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 764.365 0.070 764.435 ;
    END
  END wd_in_w1[193]
  PIN wd_in_w1[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 764.925 0.070 764.995 ;
    END
  END wd_in_w1[194]
  PIN wd_in_w1[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 765.485 0.070 765.555 ;
    END
  END wd_in_w1[195]
  PIN wd_in_w1[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 766.045 0.070 766.115 ;
    END
  END wd_in_w1[196]
  PIN wd_in_w1[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 766.605 0.070 766.675 ;
    END
  END wd_in_w1[197]
  PIN wd_in_w1[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 767.165 0.070 767.235 ;
    END
  END wd_in_w1[198]
  PIN wd_in_w1[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 767.725 0.070 767.795 ;
    END
  END wd_in_w1[199]
  PIN wd_in_w1[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 768.285 0.070 768.355 ;
    END
  END wd_in_w1[200]
  PIN wd_in_w1[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 768.845 0.070 768.915 ;
    END
  END wd_in_w1[201]
  PIN wd_in_w1[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 769.405 0.070 769.475 ;
    END
  END wd_in_w1[202]
  PIN wd_in_w1[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 769.965 0.070 770.035 ;
    END
  END wd_in_w1[203]
  PIN wd_in_w1[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 770.525 0.070 770.595 ;
    END
  END wd_in_w1[204]
  PIN wd_in_w1[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 771.085 0.070 771.155 ;
    END
  END wd_in_w1[205]
  PIN wd_in_w1[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 771.645 0.070 771.715 ;
    END
  END wd_in_w1[206]
  PIN wd_in_w1[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 772.205 0.070 772.275 ;
    END
  END wd_in_w1[207]
  PIN wd_in_w1[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 772.765 0.070 772.835 ;
    END
  END wd_in_w1[208]
  PIN wd_in_w1[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 773.325 0.070 773.395 ;
    END
  END wd_in_w1[209]
  PIN wd_in_w1[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 773.885 0.070 773.955 ;
    END
  END wd_in_w1[210]
  PIN wd_in_w1[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 774.445 0.070 774.515 ;
    END
  END wd_in_w1[211]
  PIN wd_in_w1[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 775.005 0.070 775.075 ;
    END
  END wd_in_w1[212]
  PIN wd_in_w1[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 775.565 0.070 775.635 ;
    END
  END wd_in_w1[213]
  PIN wd_in_w1[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 776.125 0.070 776.195 ;
    END
  END wd_in_w1[214]
  PIN wd_in_w1[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 776.685 0.070 776.755 ;
    END
  END wd_in_w1[215]
  PIN wd_in_w1[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 777.245 0.070 777.315 ;
    END
  END wd_in_w1[216]
  PIN wd_in_w1[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 777.805 0.070 777.875 ;
    END
  END wd_in_w1[217]
  PIN wd_in_w1[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 778.365 0.070 778.435 ;
    END
  END wd_in_w1[218]
  PIN wd_in_w1[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 778.925 0.070 778.995 ;
    END
  END wd_in_w1[219]
  PIN wd_in_w1[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 779.485 0.070 779.555 ;
    END
  END wd_in_w1[220]
  PIN wd_in_w1[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 780.045 0.070 780.115 ;
    END
  END wd_in_w1[221]
  PIN wd_in_w1[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 780.605 0.070 780.675 ;
    END
  END wd_in_w1[222]
  PIN wd_in_w1[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 781.165 0.070 781.235 ;
    END
  END wd_in_w1[223]
  PIN wd_in_w1[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 781.725 0.070 781.795 ;
    END
  END wd_in_w1[224]
  PIN wd_in_w1[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 782.285 0.070 782.355 ;
    END
  END wd_in_w1[225]
  PIN wd_in_w1[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 782.845 0.070 782.915 ;
    END
  END wd_in_w1[226]
  PIN wd_in_w1[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 783.405 0.070 783.475 ;
    END
  END wd_in_w1[227]
  PIN wd_in_w1[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 783.965 0.070 784.035 ;
    END
  END wd_in_w1[228]
  PIN wd_in_w1[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 784.525 0.070 784.595 ;
    END
  END wd_in_w1[229]
  PIN wd_in_w1[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 785.085 0.070 785.155 ;
    END
  END wd_in_w1[230]
  PIN wd_in_w1[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 785.645 0.070 785.715 ;
    END
  END wd_in_w1[231]
  PIN wd_in_w1[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 786.205 0.070 786.275 ;
    END
  END wd_in_w1[232]
  PIN wd_in_w1[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 786.765 0.070 786.835 ;
    END
  END wd_in_w1[233]
  PIN wd_in_w1[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 787.325 0.070 787.395 ;
    END
  END wd_in_w1[234]
  PIN wd_in_w1[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 787.885 0.070 787.955 ;
    END
  END wd_in_w1[235]
  PIN wd_in_w1[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 788.445 0.070 788.515 ;
    END
  END wd_in_w1[236]
  PIN wd_in_w1[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 789.005 0.070 789.075 ;
    END
  END wd_in_w1[237]
  PIN wd_in_w1[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 789.565 0.070 789.635 ;
    END
  END wd_in_w1[238]
  PIN wd_in_w1[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 790.125 0.070 790.195 ;
    END
  END wd_in_w1[239]
  PIN wd_in_w1[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 790.685 0.070 790.755 ;
    END
  END wd_in_w1[240]
  PIN wd_in_w1[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 791.245 0.070 791.315 ;
    END
  END wd_in_w1[241]
  PIN wd_in_w1[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 791.805 0.070 791.875 ;
    END
  END wd_in_w1[242]
  PIN wd_in_w1[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 792.365 0.070 792.435 ;
    END
  END wd_in_w1[243]
  PIN wd_in_w1[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 792.925 0.070 792.995 ;
    END
  END wd_in_w1[244]
  PIN wd_in_w1[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 793.485 0.070 793.555 ;
    END
  END wd_in_w1[245]
  PIN wd_in_w1[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 794.045 0.070 794.115 ;
    END
  END wd_in_w1[246]
  PIN wd_in_w1[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 794.605 0.070 794.675 ;
    END
  END wd_in_w1[247]
  PIN wd_in_w1[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 795.165 0.070 795.235 ;
    END
  END wd_in_w1[248]
  PIN wd_in_w1[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 795.725 0.070 795.795 ;
    END
  END wd_in_w1[249]
  PIN wd_in_w1[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 796.285 0.070 796.355 ;
    END
  END wd_in_w1[250]
  PIN wd_in_w1[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 796.845 0.070 796.915 ;
    END
  END wd_in_w1[251]
  PIN wd_in_w1[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 797.405 0.070 797.475 ;
    END
  END wd_in_w1[252]
  PIN wd_in_w1[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 797.965 0.070 798.035 ;
    END
  END wd_in_w1[253]
  PIN wd_in_w1[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 798.525 0.070 798.595 ;
    END
  END wd_in_w1[254]
  PIN wd_in_w1[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 799.085 0.070 799.155 ;
    END
  END wd_in_w1[255]
  PIN wd_in_w1[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 799.645 0.070 799.715 ;
    END
  END wd_in_w1[256]
  PIN wd_in_w1[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 800.205 0.070 800.275 ;
    END
  END wd_in_w1[257]
  PIN wd_in_w1[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 800.765 0.070 800.835 ;
    END
  END wd_in_w1[258]
  PIN wd_in_w1[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 801.325 0.070 801.395 ;
    END
  END wd_in_w1[259]
  PIN wd_in_w1[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 801.885 0.070 801.955 ;
    END
  END wd_in_w1[260]
  PIN wd_in_w1[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 802.445 0.070 802.515 ;
    END
  END wd_in_w1[261]
  PIN wd_in_w1[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 803.005 0.070 803.075 ;
    END
  END wd_in_w1[262]
  PIN wd_in_w1[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 803.565 0.070 803.635 ;
    END
  END wd_in_w1[263]
  PIN wd_in_w1[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 804.125 0.070 804.195 ;
    END
  END wd_in_w1[264]
  PIN wd_in_w1[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 804.685 0.070 804.755 ;
    END
  END wd_in_w1[265]
  PIN wd_in_w1[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 805.245 0.070 805.315 ;
    END
  END wd_in_w1[266]
  PIN wd_in_w1[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 805.805 0.070 805.875 ;
    END
  END wd_in_w1[267]
  PIN wd_in_w1[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 806.365 0.070 806.435 ;
    END
  END wd_in_w1[268]
  PIN wd_in_w1[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 806.925 0.070 806.995 ;
    END
  END wd_in_w1[269]
  PIN wd_in_w1[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 807.485 0.070 807.555 ;
    END
  END wd_in_w1[270]
  PIN wd_in_w1[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 808.045 0.070 808.115 ;
    END
  END wd_in_w1[271]
  PIN wd_in_w1[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 808.605 0.070 808.675 ;
    END
  END wd_in_w1[272]
  PIN wd_in_w1[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 809.165 0.070 809.235 ;
    END
  END wd_in_w1[273]
  PIN wd_in_w1[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 809.725 0.070 809.795 ;
    END
  END wd_in_w1[274]
  PIN wd_in_w1[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 810.285 0.070 810.355 ;
    END
  END wd_in_w1[275]
  PIN wd_in_w1[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 810.845 0.070 810.915 ;
    END
  END wd_in_w1[276]
  PIN wd_in_w1[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 811.405 0.070 811.475 ;
    END
  END wd_in_w1[277]
  PIN wd_in_w1[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 811.965 0.070 812.035 ;
    END
  END wd_in_w1[278]
  PIN wd_in_w1[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 812.525 0.070 812.595 ;
    END
  END wd_in_w1[279]
  PIN wd_in_w1[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 813.085 0.070 813.155 ;
    END
  END wd_in_w1[280]
  PIN wd_in_w1[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 813.645 0.070 813.715 ;
    END
  END wd_in_w1[281]
  PIN wd_in_w1[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 814.205 0.070 814.275 ;
    END
  END wd_in_w1[282]
  PIN wd_in_w1[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 814.765 0.070 814.835 ;
    END
  END wd_in_w1[283]
  PIN wd_in_w1[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 815.325 0.070 815.395 ;
    END
  END wd_in_w1[284]
  PIN wd_in_w1[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 815.885 0.070 815.955 ;
    END
  END wd_in_w1[285]
  PIN wd_in_w1[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 816.445 0.070 816.515 ;
    END
  END wd_in_w1[286]
  PIN wd_in_w1[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 817.005 0.070 817.075 ;
    END
  END wd_in_w1[287]
  PIN wd_in_w1[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 817.565 0.070 817.635 ;
    END
  END wd_in_w1[288]
  PIN wd_in_w1[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 818.125 0.070 818.195 ;
    END
  END wd_in_w1[289]
  PIN wd_in_w1[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 818.685 0.070 818.755 ;
    END
  END wd_in_w1[290]
  PIN wd_in_w1[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 819.245 0.070 819.315 ;
    END
  END wd_in_w1[291]
  PIN wd_in_w1[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 819.805 0.070 819.875 ;
    END
  END wd_in_w1[292]
  PIN wd_in_w1[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 820.365 0.070 820.435 ;
    END
  END wd_in_w1[293]
  PIN wd_in_w1[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 820.925 0.070 820.995 ;
    END
  END wd_in_w1[294]
  PIN wd_in_w1[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 821.485 0.070 821.555 ;
    END
  END wd_in_w1[295]
  PIN wd_in_w1[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 822.045 0.070 822.115 ;
    END
  END wd_in_w1[296]
  PIN wd_in_w1[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 822.605 0.070 822.675 ;
    END
  END wd_in_w1[297]
  PIN wd_in_w1[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 823.165 0.070 823.235 ;
    END
  END wd_in_w1[298]
  PIN wd_in_w1[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 823.725 0.070 823.795 ;
    END
  END wd_in_w1[299]
  PIN wd_in_w1[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 824.285 0.070 824.355 ;
    END
  END wd_in_w1[300]
  PIN wd_in_w1[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 824.845 0.070 824.915 ;
    END
  END wd_in_w1[301]
  PIN wd_in_w1[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 825.405 0.070 825.475 ;
    END
  END wd_in_w1[302]
  PIN wd_in_w1[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 825.965 0.070 826.035 ;
    END
  END wd_in_w1[303]
  PIN wd_in_w1[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 826.525 0.070 826.595 ;
    END
  END wd_in_w1[304]
  PIN wd_in_w1[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 827.085 0.070 827.155 ;
    END
  END wd_in_w1[305]
  PIN wd_in_w1[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 827.645 0.070 827.715 ;
    END
  END wd_in_w1[306]
  PIN wd_in_w1[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 828.205 0.070 828.275 ;
    END
  END wd_in_w1[307]
  PIN wd_in_w1[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 828.765 0.070 828.835 ;
    END
  END wd_in_w1[308]
  PIN wd_in_w1[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 829.325 0.070 829.395 ;
    END
  END wd_in_w1[309]
  PIN wd_in_w1[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 829.885 0.070 829.955 ;
    END
  END wd_in_w1[310]
  PIN wd_in_w1[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 830.445 0.070 830.515 ;
    END
  END wd_in_w1[311]
  PIN wd_in_w1[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.005 0.070 831.075 ;
    END
  END wd_in_w1[312]
  PIN wd_in_w1[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.565 0.070 831.635 ;
    END
  END wd_in_w1[313]
  PIN wd_in_w1[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 832.125 0.070 832.195 ;
    END
  END wd_in_w1[314]
  PIN wd_in_w1[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 832.685 0.070 832.755 ;
    END
  END wd_in_w1[315]
  PIN wd_in_w1[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 833.245 0.070 833.315 ;
    END
  END wd_in_w1[316]
  PIN wd_in_w1[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 833.805 0.070 833.875 ;
    END
  END wd_in_w1[317]
  PIN wd_in_w1[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 834.365 0.070 834.435 ;
    END
  END wd_in_w1[318]
  PIN wd_in_w1[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 834.925 0.070 834.995 ;
    END
  END wd_in_w1[319]
  PIN wd_in_w1[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 835.485 0.070 835.555 ;
    END
  END wd_in_w1[320]
  PIN wd_in_w1[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 836.045 0.070 836.115 ;
    END
  END wd_in_w1[321]
  PIN wd_in_w1[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 836.605 0.070 836.675 ;
    END
  END wd_in_w1[322]
  PIN wd_in_w1[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 837.165 0.070 837.235 ;
    END
  END wd_in_w1[323]
  PIN wd_in_w1[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 837.725 0.070 837.795 ;
    END
  END wd_in_w1[324]
  PIN wd_in_w1[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 838.285 0.070 838.355 ;
    END
  END wd_in_w1[325]
  PIN wd_in_w1[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 838.845 0.070 838.915 ;
    END
  END wd_in_w1[326]
  PIN wd_in_w1[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 839.405 0.070 839.475 ;
    END
  END wd_in_w1[327]
  PIN wd_in_w1[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 839.965 0.070 840.035 ;
    END
  END wd_in_w1[328]
  PIN wd_in_w1[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 840.525 0.070 840.595 ;
    END
  END wd_in_w1[329]
  PIN wd_in_w1[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 841.085 0.070 841.155 ;
    END
  END wd_in_w1[330]
  PIN wd_in_w1[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 841.645 0.070 841.715 ;
    END
  END wd_in_w1[331]
  PIN wd_in_w1[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 842.205 0.070 842.275 ;
    END
  END wd_in_w1[332]
  PIN wd_in_w1[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 842.765 0.070 842.835 ;
    END
  END wd_in_w1[333]
  PIN wd_in_w1[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 843.325 0.070 843.395 ;
    END
  END wd_in_w1[334]
  PIN wd_in_w1[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 843.885 0.070 843.955 ;
    END
  END wd_in_w1[335]
  PIN wd_in_w1[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 844.445 0.070 844.515 ;
    END
  END wd_in_w1[336]
  PIN wd_in_w1[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 845.005 0.070 845.075 ;
    END
  END wd_in_w1[337]
  PIN wd_in_w1[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 845.565 0.070 845.635 ;
    END
  END wd_in_w1[338]
  PIN wd_in_w1[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 846.125 0.070 846.195 ;
    END
  END wd_in_w1[339]
  PIN wd_in_w1[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 846.685 0.070 846.755 ;
    END
  END wd_in_w1[340]
  PIN wd_in_w1[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 847.245 0.070 847.315 ;
    END
  END wd_in_w1[341]
  PIN wd_in_w1[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 847.805 0.070 847.875 ;
    END
  END wd_in_w1[342]
  PIN wd_in_w1[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 848.365 0.070 848.435 ;
    END
  END wd_in_w1[343]
  PIN wd_in_w1[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 848.925 0.070 848.995 ;
    END
  END wd_in_w1[344]
  PIN wd_in_w1[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 849.485 0.070 849.555 ;
    END
  END wd_in_w1[345]
  PIN wd_in_w1[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 850.045 0.070 850.115 ;
    END
  END wd_in_w1[346]
  PIN wd_in_w1[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 850.605 0.070 850.675 ;
    END
  END wd_in_w1[347]
  PIN wd_in_w1[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 851.165 0.070 851.235 ;
    END
  END wd_in_w1[348]
  PIN wd_in_w1[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 851.725 0.070 851.795 ;
    END
  END wd_in_w1[349]
  PIN wd_in_w1[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.285 0.070 852.355 ;
    END
  END wd_in_w1[350]
  PIN wd_in_w1[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.845 0.070 852.915 ;
    END
  END wd_in_w1[351]
  PIN wd_in_w1[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 853.405 0.070 853.475 ;
    END
  END wd_in_w1[352]
  PIN wd_in_w1[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 853.965 0.070 854.035 ;
    END
  END wd_in_w1[353]
  PIN wd_in_w1[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 854.525 0.070 854.595 ;
    END
  END wd_in_w1[354]
  PIN wd_in_w1[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 855.085 0.070 855.155 ;
    END
  END wd_in_w1[355]
  PIN wd_in_w1[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 855.645 0.070 855.715 ;
    END
  END wd_in_w1[356]
  PIN wd_in_w1[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 856.205 0.070 856.275 ;
    END
  END wd_in_w1[357]
  PIN wd_in_w1[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 856.765 0.070 856.835 ;
    END
  END wd_in_w1[358]
  PIN wd_in_w1[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 857.325 0.070 857.395 ;
    END
  END wd_in_w1[359]
  PIN wd_in_w1[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 857.885 0.070 857.955 ;
    END
  END wd_in_w1[360]
  PIN wd_in_w1[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 858.445 0.070 858.515 ;
    END
  END wd_in_w1[361]
  PIN wd_in_w1[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 859.005 0.070 859.075 ;
    END
  END wd_in_w1[362]
  PIN wd_in_w1[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 859.565 0.070 859.635 ;
    END
  END wd_in_w1[363]
  PIN wd_in_w1[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 860.125 0.070 860.195 ;
    END
  END wd_in_w1[364]
  PIN wd_in_w1[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 860.685 0.070 860.755 ;
    END
  END wd_in_w1[365]
  PIN wd_in_w1[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 861.245 0.070 861.315 ;
    END
  END wd_in_w1[366]
  PIN wd_in_w1[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 861.805 0.070 861.875 ;
    END
  END wd_in_w1[367]
  PIN wd_in_w1[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 862.365 0.070 862.435 ;
    END
  END wd_in_w1[368]
  PIN wd_in_w1[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 862.925 0.070 862.995 ;
    END
  END wd_in_w1[369]
  PIN wd_in_w1[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 863.485 0.070 863.555 ;
    END
  END wd_in_w1[370]
  PIN wd_in_w1[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 864.045 0.070 864.115 ;
    END
  END wd_in_w1[371]
  PIN wd_in_w1[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 864.605 0.070 864.675 ;
    END
  END wd_in_w1[372]
  PIN wd_in_w1[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 865.165 0.070 865.235 ;
    END
  END wd_in_w1[373]
  PIN wd_in_w1[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 865.725 0.070 865.795 ;
    END
  END wd_in_w1[374]
  PIN wd_in_w1[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 866.285 0.070 866.355 ;
    END
  END wd_in_w1[375]
  PIN wd_in_w1[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 866.845 0.070 866.915 ;
    END
  END wd_in_w1[376]
  PIN wd_in_w1[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 867.405 0.070 867.475 ;
    END
  END wd_in_w1[377]
  PIN wd_in_w1[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 867.965 0.070 868.035 ;
    END
  END wd_in_w1[378]
  PIN wd_in_w1[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 868.525 0.070 868.595 ;
    END
  END wd_in_w1[379]
  PIN wd_in_w1[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 869.085 0.070 869.155 ;
    END
  END wd_in_w1[380]
  PIN wd_in_w1[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 869.645 0.070 869.715 ;
    END
  END wd_in_w1[381]
  PIN wd_in_w1[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 870.205 0.070 870.275 ;
    END
  END wd_in_w1[382]
  PIN wd_in_w1[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 870.765 0.070 870.835 ;
    END
  END wd_in_w1[383]
  PIN wd_in_w1[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 871.325 0.070 871.395 ;
    END
  END wd_in_w1[384]
  PIN wd_in_w1[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 871.885 0.070 871.955 ;
    END
  END wd_in_w1[385]
  PIN wd_in_w1[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 872.445 0.070 872.515 ;
    END
  END wd_in_w1[386]
  PIN wd_in_w1[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.005 0.070 873.075 ;
    END
  END wd_in_w1[387]
  PIN wd_in_w1[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.565 0.070 873.635 ;
    END
  END wd_in_w1[388]
  PIN wd_in_w1[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 874.125 0.070 874.195 ;
    END
  END wd_in_w1[389]
  PIN wd_in_w1[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 874.685 0.070 874.755 ;
    END
  END wd_in_w1[390]
  PIN wd_in_w1[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 875.245 0.070 875.315 ;
    END
  END wd_in_w1[391]
  PIN wd_in_w1[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 875.805 0.070 875.875 ;
    END
  END wd_in_w1[392]
  PIN wd_in_w1[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 876.365 0.070 876.435 ;
    END
  END wd_in_w1[393]
  PIN wd_in_w1[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 876.925 0.070 876.995 ;
    END
  END wd_in_w1[394]
  PIN wd_in_w1[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 877.485 0.070 877.555 ;
    END
  END wd_in_w1[395]
  PIN wd_in_w1[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 878.045 0.070 878.115 ;
    END
  END wd_in_w1[396]
  PIN wd_in_w1[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 878.605 0.070 878.675 ;
    END
  END wd_in_w1[397]
  PIN wd_in_w1[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 879.165 0.070 879.235 ;
    END
  END wd_in_w1[398]
  PIN wd_in_w1[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 879.725 0.070 879.795 ;
    END
  END wd_in_w1[399]
  PIN wd_in_w1[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 880.285 0.070 880.355 ;
    END
  END wd_in_w1[400]
  PIN wd_in_w1[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 880.845 0.070 880.915 ;
    END
  END wd_in_w1[401]
  PIN wd_in_w1[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 881.405 0.070 881.475 ;
    END
  END wd_in_w1[402]
  PIN wd_in_w1[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 881.965 0.070 882.035 ;
    END
  END wd_in_w1[403]
  PIN wd_in_w1[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 882.525 0.070 882.595 ;
    END
  END wd_in_w1[404]
  PIN wd_in_w1[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 883.085 0.070 883.155 ;
    END
  END wd_in_w1[405]
  PIN wd_in_w1[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 883.645 0.070 883.715 ;
    END
  END wd_in_w1[406]
  PIN wd_in_w1[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 884.205 0.070 884.275 ;
    END
  END wd_in_w1[407]
  PIN wd_in_w1[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 884.765 0.070 884.835 ;
    END
  END wd_in_w1[408]
  PIN wd_in_w1[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 885.325 0.070 885.395 ;
    END
  END wd_in_w1[409]
  PIN wd_in_w1[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 885.885 0.070 885.955 ;
    END
  END wd_in_w1[410]
  PIN wd_in_w1[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 886.445 0.070 886.515 ;
    END
  END wd_in_w1[411]
  PIN wd_in_w1[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 887.005 0.070 887.075 ;
    END
  END wd_in_w1[412]
  PIN wd_in_w1[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 887.565 0.070 887.635 ;
    END
  END wd_in_w1[413]
  PIN wd_in_w1[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 888.125 0.070 888.195 ;
    END
  END wd_in_w1[414]
  PIN wd_in_w1[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 888.685 0.070 888.755 ;
    END
  END wd_in_w1[415]
  PIN wd_in_w1[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 889.245 0.070 889.315 ;
    END
  END wd_in_w1[416]
  PIN wd_in_w1[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 889.805 0.070 889.875 ;
    END
  END wd_in_w1[417]
  PIN wd_in_w1[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 890.365 0.070 890.435 ;
    END
  END wd_in_w1[418]
  PIN wd_in_w1[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 890.925 0.070 890.995 ;
    END
  END wd_in_w1[419]
  PIN wd_in_w1[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 891.485 0.070 891.555 ;
    END
  END wd_in_w1[420]
  PIN wd_in_w1[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 892.045 0.070 892.115 ;
    END
  END wd_in_w1[421]
  PIN wd_in_w1[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 892.605 0.070 892.675 ;
    END
  END wd_in_w1[422]
  PIN wd_in_w1[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 893.165 0.070 893.235 ;
    END
  END wd_in_w1[423]
  PIN wd_in_w1[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 893.725 0.070 893.795 ;
    END
  END wd_in_w1[424]
  PIN wd_in_w1[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 894.285 0.070 894.355 ;
    END
  END wd_in_w1[425]
  PIN wd_in_w1[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 894.845 0.070 894.915 ;
    END
  END wd_in_w1[426]
  PIN wd_in_w1[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 895.405 0.070 895.475 ;
    END
  END wd_in_w1[427]
  PIN wd_in_w1[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 895.965 0.070 896.035 ;
    END
  END wd_in_w1[428]
  PIN wd_in_w1[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 896.525 0.070 896.595 ;
    END
  END wd_in_w1[429]
  PIN wd_in_w1[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 897.085 0.070 897.155 ;
    END
  END wd_in_w1[430]
  PIN wd_in_w1[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 897.645 0.070 897.715 ;
    END
  END wd_in_w1[431]
  PIN wd_in_w1[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 898.205 0.070 898.275 ;
    END
  END wd_in_w1[432]
  PIN wd_in_w1[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 898.765 0.070 898.835 ;
    END
  END wd_in_w1[433]
  PIN wd_in_w1[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 899.325 0.070 899.395 ;
    END
  END wd_in_w1[434]
  PIN wd_in_w1[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 899.885 0.070 899.955 ;
    END
  END wd_in_w1[435]
  PIN wd_in_w1[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 900.445 0.070 900.515 ;
    END
  END wd_in_w1[436]
  PIN wd_in_w1[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 901.005 0.070 901.075 ;
    END
  END wd_in_w1[437]
  PIN wd_in_w1[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 901.565 0.070 901.635 ;
    END
  END wd_in_w1[438]
  PIN wd_in_w1[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 902.125 0.070 902.195 ;
    END
  END wd_in_w1[439]
  PIN wd_in_w1[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 902.685 0.070 902.755 ;
    END
  END wd_in_w1[440]
  PIN wd_in_w1[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 903.245 0.070 903.315 ;
    END
  END wd_in_w1[441]
  PIN wd_in_w1[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 903.805 0.070 903.875 ;
    END
  END wd_in_w1[442]
  PIN wd_in_w1[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 904.365 0.070 904.435 ;
    END
  END wd_in_w1[443]
  PIN wd_in_w1[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 904.925 0.070 904.995 ;
    END
  END wd_in_w1[444]
  PIN wd_in_w1[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 905.485 0.070 905.555 ;
    END
  END wd_in_w1[445]
  PIN wd_in_w1[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 906.045 0.070 906.115 ;
    END
  END wd_in_w1[446]
  PIN wd_in_w1[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 906.605 0.070 906.675 ;
    END
  END wd_in_w1[447]
  PIN wd_in_w1[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 907.165 0.070 907.235 ;
    END
  END wd_in_w1[448]
  PIN wd_in_w1[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 907.725 0.070 907.795 ;
    END
  END wd_in_w1[449]
  PIN wd_in_w1[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 908.285 0.070 908.355 ;
    END
  END wd_in_w1[450]
  PIN wd_in_w1[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 908.845 0.070 908.915 ;
    END
  END wd_in_w1[451]
  PIN wd_in_w1[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 909.405 0.070 909.475 ;
    END
  END wd_in_w1[452]
  PIN wd_in_w1[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 909.965 0.070 910.035 ;
    END
  END wd_in_w1[453]
  PIN wd_in_w1[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 910.525 0.070 910.595 ;
    END
  END wd_in_w1[454]
  PIN wd_in_w1[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 911.085 0.070 911.155 ;
    END
  END wd_in_w1[455]
  PIN wd_in_w1[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 911.645 0.070 911.715 ;
    END
  END wd_in_w1[456]
  PIN wd_in_w1[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 912.205 0.070 912.275 ;
    END
  END wd_in_w1[457]
  PIN wd_in_w1[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 912.765 0.070 912.835 ;
    END
  END wd_in_w1[458]
  PIN wd_in_w1[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 913.325 0.070 913.395 ;
    END
  END wd_in_w1[459]
  PIN wd_in_w1[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 913.885 0.070 913.955 ;
    END
  END wd_in_w1[460]
  PIN wd_in_w1[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 914.445 0.070 914.515 ;
    END
  END wd_in_w1[461]
  PIN wd_in_w1[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 915.005 0.070 915.075 ;
    END
  END wd_in_w1[462]
  PIN wd_in_w1[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 915.565 0.070 915.635 ;
    END
  END wd_in_w1[463]
  PIN wd_in_w1[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 916.125 0.070 916.195 ;
    END
  END wd_in_w1[464]
  PIN wd_in_w1[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 916.685 0.070 916.755 ;
    END
  END wd_in_w1[465]
  PIN wd_in_w1[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 917.245 0.070 917.315 ;
    END
  END wd_in_w1[466]
  PIN wd_in_w1[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 917.805 0.070 917.875 ;
    END
  END wd_in_w1[467]
  PIN wd_in_w1[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 918.365 0.070 918.435 ;
    END
  END wd_in_w1[468]
  PIN wd_in_w1[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 918.925 0.070 918.995 ;
    END
  END wd_in_w1[469]
  PIN wd_in_w1[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 919.485 0.070 919.555 ;
    END
  END wd_in_w1[470]
  PIN wd_in_w1[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 920.045 0.070 920.115 ;
    END
  END wd_in_w1[471]
  PIN wd_in_w1[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 920.605 0.070 920.675 ;
    END
  END wd_in_w1[472]
  PIN wd_in_w1[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 921.165 0.070 921.235 ;
    END
  END wd_in_w1[473]
  PIN wd_in_w1[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 921.725 0.070 921.795 ;
    END
  END wd_in_w1[474]
  PIN wd_in_w1[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 922.285 0.070 922.355 ;
    END
  END wd_in_w1[475]
  PIN wd_in_w1[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 922.845 0.070 922.915 ;
    END
  END wd_in_w1[476]
  PIN wd_in_w1[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 923.405 0.070 923.475 ;
    END
  END wd_in_w1[477]
  PIN wd_in_w1[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 923.965 0.070 924.035 ;
    END
  END wd_in_w1[478]
  PIN wd_in_w1[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 924.525 0.070 924.595 ;
    END
  END wd_in_w1[479]
  PIN wd_in_w1[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 925.085 0.070 925.155 ;
    END
  END wd_in_w1[480]
  PIN wd_in_w1[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 925.645 0.070 925.715 ;
    END
  END wd_in_w1[481]
  PIN wd_in_w1[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 926.205 0.070 926.275 ;
    END
  END wd_in_w1[482]
  PIN wd_in_w1[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 926.765 0.070 926.835 ;
    END
  END wd_in_w1[483]
  PIN wd_in_w1[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 927.325 0.070 927.395 ;
    END
  END wd_in_w1[484]
  PIN wd_in_w1[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 927.885 0.070 927.955 ;
    END
  END wd_in_w1[485]
  PIN wd_in_w1[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 928.445 0.070 928.515 ;
    END
  END wd_in_w1[486]
  PIN wd_in_w1[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 929.005 0.070 929.075 ;
    END
  END wd_in_w1[487]
  PIN wd_in_w1[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 929.565 0.070 929.635 ;
    END
  END wd_in_w1[488]
  PIN wd_in_w1[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 930.125 0.070 930.195 ;
    END
  END wd_in_w1[489]
  PIN wd_in_w1[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 930.685 0.070 930.755 ;
    END
  END wd_in_w1[490]
  PIN wd_in_w1[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 931.245 0.070 931.315 ;
    END
  END wd_in_w1[491]
  PIN wd_in_w1[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 931.805 0.070 931.875 ;
    END
  END wd_in_w1[492]
  PIN wd_in_w1[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 932.365 0.070 932.435 ;
    END
  END wd_in_w1[493]
  PIN wd_in_w1[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 932.925 0.070 932.995 ;
    END
  END wd_in_w1[494]
  PIN wd_in_w1[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 933.485 0.070 933.555 ;
    END
  END wd_in_w1[495]
  PIN wd_in_w1[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 934.045 0.070 934.115 ;
    END
  END wd_in_w1[496]
  PIN wd_in_w1[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 934.605 0.070 934.675 ;
    END
  END wd_in_w1[497]
  PIN wd_in_w1[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 935.165 0.070 935.235 ;
    END
  END wd_in_w1[498]
  PIN wd_in_w1[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 935.725 0.070 935.795 ;
    END
  END wd_in_w1[499]
  PIN wd_in_w1[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 936.285 0.070 936.355 ;
    END
  END wd_in_w1[500]
  PIN wd_in_w1[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 936.845 0.070 936.915 ;
    END
  END wd_in_w1[501]
  PIN wd_in_w1[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 937.405 0.070 937.475 ;
    END
  END wd_in_w1[502]
  PIN wd_in_w1[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 937.965 0.070 938.035 ;
    END
  END wd_in_w1[503]
  PIN wd_in_w1[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 938.525 0.070 938.595 ;
    END
  END wd_in_w1[504]
  PIN wd_in_w1[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 939.085 0.070 939.155 ;
    END
  END wd_in_w1[505]
  PIN wd_in_w1[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 939.645 0.070 939.715 ;
    END
  END wd_in_w1[506]
  PIN wd_in_w1[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 940.205 0.070 940.275 ;
    END
  END wd_in_w1[507]
  PIN wd_in_w1[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 940.765 0.070 940.835 ;
    END
  END wd_in_w1[508]
  PIN wd_in_w1[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 941.325 0.070 941.395 ;
    END
  END wd_in_w1[509]
  PIN wd_in_w1[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 941.885 0.070 941.955 ;
    END
  END wd_in_w1[510]
  PIN wd_in_w1[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 942.445 0.070 942.515 ;
    END
  END wd_in_w1[511]
  PIN addr_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 970.165 0.070 970.235 ;
    END
  END addr_w1[0]
  PIN addr_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 970.725 0.070 970.795 ;
    END
  END addr_w1[1]
  PIN addr_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 971.285 0.070 971.355 ;
    END
  END addr_w1[2]
  PIN addr_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 971.845 0.070 971.915 ;
    END
  END addr_w1[3]
  PIN addr_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 972.405 0.070 972.475 ;
    END
  END addr_w1[4]
  PIN addr_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 972.965 0.070 973.035 ;
    END
  END addr_w1[5]
  PIN addr_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 973.525 0.070 973.595 ;
    END
  END addr_w1[6]
  PIN addr_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 974.085 0.070 974.155 ;
    END
  END addr_w1[7]
  PIN addr_w1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 974.645 0.070 974.715 ;
    END
  END addr_w1[8]
  PIN addr_w1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 975.205 0.070 975.275 ;
    END
  END addr_w1[9]
  PIN addr_r1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1002.925 0.070 1002.995 ;
    END
  END addr_r1[0]
  PIN addr_r1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1003.485 0.070 1003.555 ;
    END
  END addr_r1[1]
  PIN addr_r1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1004.045 0.070 1004.115 ;
    END
  END addr_r1[2]
  PIN addr_r1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1004.605 0.070 1004.675 ;
    END
  END addr_r1[3]
  PIN addr_r1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1005.165 0.070 1005.235 ;
    END
  END addr_r1[4]
  PIN addr_r1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1005.725 0.070 1005.795 ;
    END
  END addr_r1[5]
  PIN addr_r1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1006.285 0.070 1006.355 ;
    END
  END addr_r1[6]
  PIN addr_r1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1006.845 0.070 1006.915 ;
    END
  END addr_r1[7]
  PIN addr_r1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1007.405 0.070 1007.475 ;
    END
  END addr_r1[8]
  PIN addr_r1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1007.965 0.070 1008.035 ;
    END
  END addr_r1[9]
  PIN we_in_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1035.685 0.070 1035.755 ;
    END
  END we_in_w1
  PIN ce_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1090.565 0.070 1090.635 ;
    END
  END ce_w1
  PIN ce_r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1118.285 0.070 1118.355 ;
    END
  END ce_r1
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1146.005 0.070 1146.075 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 980.000 ;
      RECT 3.500 1.400 3.780 980.000 ;
      RECT 5.740 1.400 6.020 980.000 ;
      RECT 7.980 1.400 8.260 980.000 ;
      RECT 10.220 1.400 10.500 980.000 ;
      RECT 12.460 1.400 12.740 980.000 ;
      RECT 14.700 1.400 14.980 980.000 ;
      RECT 16.940 1.400 17.220 980.000 ;
      RECT 19.180 1.400 19.460 980.000 ;
      RECT 21.420 1.400 21.700 980.000 ;
      RECT 23.660 1.400 23.940 980.000 ;
      RECT 25.900 1.400 26.180 980.000 ;
      RECT 28.140 1.400 28.420 980.000 ;
      RECT 30.380 1.400 30.660 980.000 ;
      RECT 32.620 1.400 32.900 980.000 ;
      RECT 34.860 1.400 35.140 980.000 ;
      RECT 37.100 1.400 37.380 980.000 ;
      RECT 39.340 1.400 39.620 980.000 ;
      RECT 41.580 1.400 41.860 980.000 ;
      RECT 43.820 1.400 44.100 980.000 ;
      RECT 46.060 1.400 46.340 980.000 ;
      RECT 48.300 1.400 48.580 980.000 ;
      RECT 50.540 1.400 50.820 980.000 ;
      RECT 52.780 1.400 53.060 980.000 ;
      RECT 55.020 1.400 55.300 980.000 ;
      RECT 57.260 1.400 57.540 980.000 ;
      RECT 59.500 1.400 59.780 980.000 ;
      RECT 61.740 1.400 62.020 980.000 ;
      RECT 63.980 1.400 64.260 980.000 ;
      RECT 66.220 1.400 66.500 980.000 ;
      RECT 68.460 1.400 68.740 980.000 ;
      RECT 70.700 1.400 70.980 980.000 ;
      RECT 72.940 1.400 73.220 980.000 ;
      RECT 75.180 1.400 75.460 980.000 ;
      RECT 77.420 1.400 77.700 980.000 ;
      RECT 79.660 1.400 79.940 980.000 ;
      RECT 81.900 1.400 82.180 980.000 ;
      RECT 84.140 1.400 84.420 980.000 ;
      RECT 86.380 1.400 86.660 980.000 ;
      RECT 88.620 1.400 88.900 980.000 ;
      RECT 90.860 1.400 91.140 980.000 ;
      RECT 93.100 1.400 93.380 980.000 ;
      RECT 95.340 1.400 95.620 980.000 ;
      RECT 97.580 1.400 97.860 980.000 ;
      RECT 99.820 1.400 100.100 980.000 ;
      RECT 102.060 1.400 102.340 980.000 ;
      RECT 104.300 1.400 104.580 980.000 ;
      RECT 106.540 1.400 106.820 980.000 ;
      RECT 108.780 1.400 109.060 980.000 ;
      RECT 111.020 1.400 111.300 980.000 ;
      RECT 113.260 1.400 113.540 980.000 ;
      RECT 115.500 1.400 115.780 980.000 ;
      RECT 117.740 1.400 118.020 980.000 ;
      RECT 119.980 1.400 120.260 980.000 ;
      RECT 122.220 1.400 122.500 980.000 ;
      RECT 124.460 1.400 124.740 980.000 ;
      RECT 126.700 1.400 126.980 980.000 ;
      RECT 128.940 1.400 129.220 980.000 ;
      RECT 131.180 1.400 131.460 980.000 ;
      RECT 133.420 1.400 133.700 980.000 ;
      RECT 135.660 1.400 135.940 980.000 ;
      RECT 137.900 1.400 138.180 980.000 ;
      RECT 140.140 1.400 140.420 980.000 ;
      RECT 142.380 1.400 142.660 980.000 ;
      RECT 144.620 1.400 144.900 980.000 ;
      RECT 146.860 1.400 147.140 980.000 ;
      RECT 149.100 1.400 149.380 980.000 ;
      RECT 151.340 1.400 151.620 980.000 ;
      RECT 153.580 1.400 153.860 980.000 ;
      RECT 155.820 1.400 156.100 980.000 ;
      RECT 158.060 1.400 158.340 980.000 ;
      RECT 160.300 1.400 160.580 980.000 ;
      RECT 162.540 1.400 162.820 980.000 ;
      RECT 164.780 1.400 165.060 980.000 ;
      RECT 167.020 1.400 167.300 980.000 ;
      RECT 169.260 1.400 169.540 980.000 ;
      RECT 171.500 1.400 171.780 980.000 ;
      RECT 173.740 1.400 174.020 980.000 ;
      RECT 175.980 1.400 176.260 980.000 ;
      RECT 178.220 1.400 178.500 980.000 ;
      RECT 180.460 1.400 180.740 980.000 ;
      RECT 182.700 1.400 182.980 980.000 ;
      RECT 184.940 1.400 185.220 980.000 ;
      RECT 187.180 1.400 187.460 980.000 ;
      RECT 189.420 1.400 189.700 980.000 ;
      RECT 191.660 1.400 191.940 980.000 ;
      RECT 193.900 1.400 194.180 980.000 ;
      RECT 196.140 1.400 196.420 980.000 ;
      RECT 198.380 1.400 198.660 980.000 ;
      RECT 200.620 1.400 200.900 980.000 ;
      RECT 202.860 1.400 203.140 980.000 ;
      RECT 205.100 1.400 205.380 980.000 ;
      RECT 207.340 1.400 207.620 980.000 ;
      RECT 209.580 1.400 209.860 980.000 ;
      RECT 211.820 1.400 212.100 980.000 ;
      RECT 214.060 1.400 214.340 980.000 ;
      RECT 216.300 1.400 216.580 980.000 ;
      RECT 218.540 1.400 218.820 980.000 ;
      RECT 220.780 1.400 221.060 980.000 ;
      RECT 223.020 1.400 223.300 980.000 ;
      RECT 225.260 1.400 225.540 980.000 ;
      RECT 227.500 1.400 227.780 980.000 ;
      RECT 229.740 1.400 230.020 980.000 ;
      RECT 231.980 1.400 232.260 980.000 ;
      RECT 234.220 1.400 234.500 980.000 ;
      RECT 236.460 1.400 236.740 980.000 ;
      RECT 238.700 1.400 238.980 980.000 ;
      RECT 240.940 1.400 241.220 980.000 ;
      RECT 243.180 1.400 243.460 980.000 ;
      RECT 245.420 1.400 245.700 980.000 ;
      RECT 247.660 1.400 247.940 980.000 ;
      RECT 249.900 1.400 250.180 980.000 ;
      RECT 252.140 1.400 252.420 980.000 ;
      RECT 254.380 1.400 254.660 980.000 ;
      RECT 256.620 1.400 256.900 980.000 ;
      RECT 258.860 1.400 259.140 980.000 ;
      RECT 261.100 1.400 261.380 980.000 ;
      RECT 263.340 1.400 263.620 980.000 ;
      RECT 265.580 1.400 265.860 980.000 ;
      RECT 267.820 1.400 268.100 980.000 ;
      RECT 270.060 1.400 270.340 980.000 ;
      RECT 272.300 1.400 272.580 980.000 ;
      RECT 274.540 1.400 274.820 980.000 ;
      RECT 276.780 1.400 277.060 980.000 ;
      RECT 279.020 1.400 279.300 980.000 ;
      RECT 281.260 1.400 281.540 980.000 ;
      RECT 283.500 1.400 283.780 980.000 ;
      RECT 285.740 1.400 286.020 980.000 ;
      RECT 287.980 1.400 288.260 980.000 ;
      RECT 290.220 1.400 290.500 980.000 ;
      RECT 292.460 1.400 292.740 980.000 ;
      RECT 294.700 1.400 294.980 980.000 ;
      RECT 296.940 1.400 297.220 980.000 ;
      RECT 299.180 1.400 299.460 980.000 ;
      RECT 301.420 1.400 301.700 980.000 ;
      RECT 303.660 1.400 303.940 980.000 ;
      RECT 305.900 1.400 306.180 980.000 ;
      RECT 308.140 1.400 308.420 980.000 ;
      RECT 310.380 1.400 310.660 980.000 ;
      RECT 312.620 1.400 312.900 980.000 ;
      RECT 314.860 1.400 315.140 980.000 ;
      RECT 317.100 1.400 317.380 980.000 ;
      RECT 319.340 1.400 319.620 980.000 ;
      RECT 321.580 1.400 321.860 980.000 ;
      RECT 323.820 1.400 324.100 980.000 ;
      RECT 326.060 1.400 326.340 980.000 ;
      RECT 328.300 1.400 328.580 980.000 ;
      RECT 330.540 1.400 330.820 980.000 ;
      RECT 332.780 1.400 333.060 980.000 ;
      RECT 335.020 1.400 335.300 980.000 ;
      RECT 337.260 1.400 337.540 980.000 ;
      RECT 339.500 1.400 339.780 980.000 ;
      RECT 341.740 1.400 342.020 980.000 ;
      RECT 343.980 1.400 344.260 980.000 ;
      RECT 346.220 1.400 346.500 980.000 ;
      RECT 348.460 1.400 348.740 980.000 ;
      RECT 350.700 1.400 350.980 980.000 ;
      RECT 352.940 1.400 353.220 980.000 ;
      RECT 355.180 1.400 355.460 980.000 ;
      RECT 357.420 1.400 357.700 980.000 ;
      RECT 359.660 1.400 359.940 980.000 ;
      RECT 361.900 1.400 362.180 980.000 ;
      RECT 364.140 1.400 364.420 980.000 ;
      RECT 366.380 1.400 366.660 980.000 ;
      RECT 368.620 1.400 368.900 980.000 ;
      RECT 370.860 1.400 371.140 980.000 ;
      RECT 373.100 1.400 373.380 980.000 ;
      RECT 375.340 1.400 375.620 980.000 ;
      RECT 377.580 1.400 377.860 980.000 ;
      RECT 379.820 1.400 380.100 980.000 ;
      RECT 382.060 1.400 382.340 980.000 ;
      RECT 384.300 1.400 384.580 980.000 ;
      RECT 386.540 1.400 386.820 980.000 ;
      RECT 388.780 1.400 389.060 980.000 ;
      RECT 391.020 1.400 391.300 980.000 ;
      RECT 393.260 1.400 393.540 980.000 ;
      RECT 395.500 1.400 395.780 980.000 ;
      RECT 397.740 1.400 398.020 980.000 ;
      RECT 399.980 1.400 400.260 980.000 ;
      RECT 402.220 1.400 402.500 980.000 ;
      RECT 404.460 1.400 404.740 980.000 ;
      RECT 406.700 1.400 406.980 980.000 ;
      RECT 408.940 1.400 409.220 980.000 ;
      RECT 411.180 1.400 411.460 980.000 ;
      RECT 413.420 1.400 413.700 980.000 ;
      RECT 415.660 1.400 415.940 980.000 ;
      RECT 417.900 1.400 418.180 980.000 ;
      RECT 420.140 1.400 420.420 980.000 ;
      RECT 422.380 1.400 422.660 980.000 ;
      RECT 424.620 1.400 424.900 980.000 ;
      RECT 426.860 1.400 427.140 980.000 ;
      RECT 429.100 1.400 429.380 980.000 ;
      RECT 431.340 1.400 431.620 980.000 ;
      RECT 433.580 1.400 433.860 980.000 ;
      RECT 435.820 1.400 436.100 980.000 ;
      RECT 438.060 1.400 438.340 980.000 ;
      RECT 440.300 1.400 440.580 980.000 ;
      RECT 442.540 1.400 442.820 980.000 ;
      RECT 444.780 1.400 445.060 980.000 ;
      RECT 447.020 1.400 447.300 980.000 ;
      RECT 449.260 1.400 449.540 980.000 ;
      RECT 451.500 1.400 451.780 980.000 ;
      RECT 453.740 1.400 454.020 980.000 ;
      RECT 455.980 1.400 456.260 980.000 ;
      RECT 458.220 1.400 458.500 980.000 ;
      RECT 460.460 1.400 460.740 980.000 ;
      RECT 462.700 1.400 462.980 980.000 ;
      RECT 464.940 1.400 465.220 980.000 ;
      RECT 467.180 1.400 467.460 980.000 ;
      RECT 469.420 1.400 469.700 980.000 ;
      RECT 471.660 1.400 471.940 980.000 ;
      RECT 473.900 1.400 474.180 980.000 ;
      RECT 476.140 1.400 476.420 980.000 ;
      RECT 478.380 1.400 478.660 980.000 ;
      RECT 480.620 1.400 480.900 980.000 ;
      RECT 482.860 1.400 483.140 980.000 ;
      RECT 485.100 1.400 485.380 980.000 ;
      RECT 487.340 1.400 487.620 980.000 ;
      RECT 489.580 1.400 489.860 980.000 ;
      RECT 491.820 1.400 492.100 980.000 ;
      RECT 494.060 1.400 494.340 980.000 ;
      RECT 496.300 1.400 496.580 980.000 ;
      RECT 498.540 1.400 498.820 980.000 ;
      RECT 500.780 1.400 501.060 980.000 ;
      RECT 503.020 1.400 503.300 980.000 ;
      RECT 505.260 1.400 505.540 980.000 ;
      RECT 507.500 1.400 507.780 980.000 ;
      RECT 509.740 1.400 510.020 980.000 ;
      RECT 511.980 1.400 512.260 980.000 ;
      RECT 514.220 1.400 514.500 980.000 ;
      RECT 516.460 1.400 516.740 980.000 ;
      RECT 518.700 1.400 518.980 980.000 ;
      RECT 520.940 1.400 521.220 980.000 ;
      RECT 523.180 1.400 523.460 980.000 ;
      RECT 525.420 1.400 525.700 980.000 ;
      RECT 527.660 1.400 527.940 980.000 ;
      RECT 529.900 1.400 530.180 980.000 ;
      RECT 532.140 1.400 532.420 980.000 ;
      RECT 534.380 1.400 534.660 980.000 ;
      RECT 536.620 1.400 536.900 980.000 ;
      RECT 538.860 1.400 539.140 980.000 ;
      RECT 541.100 1.400 541.380 980.000 ;
      RECT 543.340 1.400 543.620 980.000 ;
      RECT 545.580 1.400 545.860 980.000 ;
      RECT 547.820 1.400 548.100 980.000 ;
      RECT 550.060 1.400 550.340 980.000 ;
      RECT 552.300 1.400 552.580 980.000 ;
      RECT 554.540 1.400 554.820 980.000 ;
      RECT 556.780 1.400 557.060 980.000 ;
      RECT 559.020 1.400 559.300 980.000 ;
      RECT 561.260 1.400 561.540 980.000 ;
      RECT 563.500 1.400 563.780 980.000 ;
      RECT 565.740 1.400 566.020 980.000 ;
      RECT 567.980 1.400 568.260 980.000 ;
      RECT 570.220 1.400 570.500 980.000 ;
      RECT 572.460 1.400 572.740 980.000 ;
      RECT 574.700 1.400 574.980 980.000 ;
      RECT 576.940 1.400 577.220 980.000 ;
      RECT 579.180 1.400 579.460 980.000 ;
      RECT 581.420 1.400 581.700 980.000 ;
      RECT 583.660 1.400 583.940 980.000 ;
      RECT 585.900 1.400 586.180 980.000 ;
      RECT 588.140 1.400 588.420 980.000 ;
      RECT 590.380 1.400 590.660 980.000 ;
      RECT 592.620 1.400 592.900 980.000 ;
      RECT 594.860 1.400 595.140 980.000 ;
      RECT 597.100 1.400 597.380 980.000 ;
      RECT 599.340 1.400 599.620 980.000 ;
      RECT 601.580 1.400 601.860 980.000 ;
      RECT 603.820 1.400 604.100 980.000 ;
      RECT 606.060 1.400 606.340 980.000 ;
      RECT 608.300 1.400 608.580 980.000 ;
      RECT 610.540 1.400 610.820 980.000 ;
      RECT 612.780 1.400 613.060 980.000 ;
      RECT 615.020 1.400 615.300 980.000 ;
      RECT 617.260 1.400 617.540 980.000 ;
      RECT 619.500 1.400 619.780 980.000 ;
      RECT 621.740 1.400 622.020 980.000 ;
      RECT 623.980 1.400 624.260 980.000 ;
      RECT 626.220 1.400 626.500 980.000 ;
      RECT 628.460 1.400 628.740 980.000 ;
      RECT 630.700 1.400 630.980 980.000 ;
      RECT 632.940 1.400 633.220 980.000 ;
      RECT 635.180 1.400 635.460 980.000 ;
      RECT 637.420 1.400 637.700 980.000 ;
      RECT 639.660 1.400 639.940 980.000 ;
      RECT 641.900 1.400 642.180 980.000 ;
      RECT 644.140 1.400 644.420 980.000 ;
      RECT 646.380 1.400 646.660 980.000 ;
      RECT 648.620 1.400 648.900 980.000 ;
      RECT 650.860 1.400 651.140 980.000 ;
      RECT 653.100 1.400 653.380 980.000 ;
      RECT 655.340 1.400 655.620 980.000 ;
      RECT 657.580 1.400 657.860 980.000 ;
      RECT 659.820 1.400 660.100 980.000 ;
      RECT 662.060 1.400 662.340 980.000 ;
      RECT 664.300 1.400 664.580 980.000 ;
      RECT 666.540 1.400 666.820 980.000 ;
      RECT 668.780 1.400 669.060 980.000 ;
      RECT 671.020 1.400 671.300 980.000 ;
      RECT 673.260 1.400 673.540 980.000 ;
      RECT 675.500 1.400 675.780 980.000 ;
      RECT 677.740 1.400 678.020 980.000 ;
      RECT 679.980 1.400 680.260 980.000 ;
      RECT 682.220 1.400 682.500 980.000 ;
      RECT 684.460 1.400 684.740 980.000 ;
      RECT 686.700 1.400 686.980 980.000 ;
      RECT 688.940 1.400 689.220 980.000 ;
      RECT 691.180 1.400 691.460 980.000 ;
      RECT 693.420 1.400 693.700 980.000 ;
      RECT 695.660 1.400 695.940 980.000 ;
      RECT 697.900 1.400 698.180 980.000 ;
      RECT 700.140 1.400 700.420 980.000 ;
      RECT 702.380 1.400 702.660 980.000 ;
      RECT 704.620 1.400 704.900 980.000 ;
      RECT 706.860 1.400 707.140 980.000 ;
      RECT 709.100 1.400 709.380 980.000 ;
      RECT 711.340 1.400 711.620 980.000 ;
      RECT 713.580 1.400 713.860 980.000 ;
      RECT 715.820 1.400 716.100 980.000 ;
      RECT 718.060 1.400 718.340 980.000 ;
      RECT 720.300 1.400 720.580 980.000 ;
      RECT 722.540 1.400 722.820 980.000 ;
      RECT 724.780 1.400 725.060 980.000 ;
      RECT 727.020 1.400 727.300 980.000 ;
      RECT 729.260 1.400 729.540 980.000 ;
      RECT 731.500 1.400 731.780 980.000 ;
      RECT 733.740 1.400 734.020 980.000 ;
      RECT 735.980 1.400 736.260 980.000 ;
      RECT 738.220 1.400 738.500 980.000 ;
      RECT 740.460 1.400 740.740 980.000 ;
      RECT 742.700 1.400 742.980 980.000 ;
      RECT 744.940 1.400 745.220 980.000 ;
      RECT 747.180 1.400 747.460 980.000 ;
      RECT 749.420 1.400 749.700 980.000 ;
      RECT 751.660 1.400 751.940 980.000 ;
      RECT 753.900 1.400 754.180 980.000 ;
      RECT 756.140 1.400 756.420 980.000 ;
      RECT 758.380 1.400 758.660 980.000 ;
      RECT 760.620 1.400 760.900 980.000 ;
      RECT 762.860 1.400 763.140 980.000 ;
      RECT 765.100 1.400 765.380 980.000 ;
      RECT 767.340 1.400 767.620 980.000 ;
      RECT 769.580 1.400 769.860 980.000 ;
      RECT 771.820 1.400 772.100 980.000 ;
      RECT 774.060 1.400 774.340 980.000 ;
      RECT 776.300 1.400 776.580 980.000 ;
      RECT 778.540 1.400 778.820 980.000 ;
      RECT 780.780 1.400 781.060 980.000 ;
      RECT 783.020 1.400 783.300 980.000 ;
      RECT 785.260 1.400 785.540 980.000 ;
      RECT 787.500 1.400 787.780 980.000 ;
      RECT 789.740 1.400 790.020 980.000 ;
      RECT 791.980 1.400 792.260 980.000 ;
      RECT 794.220 1.400 794.500 980.000 ;
      RECT 796.460 1.400 796.740 980.000 ;
      RECT 798.700 1.400 798.980 980.000 ;
      RECT 800.940 1.400 801.220 980.000 ;
      RECT 803.180 1.400 803.460 980.000 ;
      RECT 805.420 1.400 805.700 980.000 ;
      RECT 807.660 1.400 807.940 980.000 ;
      RECT 809.900 1.400 810.180 980.000 ;
      RECT 812.140 1.400 812.420 980.000 ;
      RECT 814.380 1.400 814.660 980.000 ;
      RECT 816.620 1.400 816.900 980.000 ;
      RECT 818.860 1.400 819.140 980.000 ;
      RECT 821.100 1.400 821.380 980.000 ;
      RECT 823.340 1.400 823.620 980.000 ;
      RECT 825.580 1.400 825.860 980.000 ;
      RECT 827.820 1.400 828.100 980.000 ;
      RECT 830.060 1.400 830.340 980.000 ;
      RECT 832.300 1.400 832.580 980.000 ;
      RECT 834.540 1.400 834.820 980.000 ;
      RECT 836.780 1.400 837.060 980.000 ;
      RECT 839.020 1.400 839.300 980.000 ;
      RECT 841.260 1.400 841.540 980.000 ;
      RECT 843.500 1.400 843.780 980.000 ;
      RECT 845.740 1.400 846.020 980.000 ;
      RECT 847.980 1.400 848.260 980.000 ;
      RECT 850.220 1.400 850.500 980.000 ;
      RECT 852.460 1.400 852.740 980.000 ;
      RECT 854.700 1.400 854.980 980.000 ;
      RECT 856.940 1.400 857.220 980.000 ;
      RECT 859.180 1.400 859.460 980.000 ;
      RECT 861.420 1.400 861.700 980.000 ;
      RECT 863.660 1.400 863.940 980.000 ;
      RECT 865.900 1.400 866.180 980.000 ;
      RECT 868.140 1.400 868.420 980.000 ;
      RECT 870.380 1.400 870.660 980.000 ;
      RECT 872.620 1.400 872.900 980.000 ;
      RECT 874.860 1.400 875.140 980.000 ;
      RECT 877.100 1.400 877.380 980.000 ;
      RECT 879.340 1.400 879.620 980.000 ;
      RECT 881.580 1.400 881.860 980.000 ;
      RECT 883.820 1.400 884.100 980.000 ;
      RECT 886.060 1.400 886.340 980.000 ;
      RECT 888.300 1.400 888.580 980.000 ;
      RECT 890.540 1.400 890.820 980.000 ;
      RECT 892.780 1.400 893.060 980.000 ;
      RECT 895.020 1.400 895.300 980.000 ;
      RECT 897.260 1.400 897.540 980.000 ;
      RECT 899.500 1.400 899.780 980.000 ;
      RECT 901.740 1.400 902.020 980.000 ;
      RECT 903.980 1.400 904.260 980.000 ;
      RECT 906.220 1.400 906.500 980.000 ;
      RECT 908.460 1.400 908.740 980.000 ;
      RECT 910.700 1.400 910.980 980.000 ;
      RECT 912.940 1.400 913.220 980.000 ;
      RECT 915.180 1.400 915.460 980.000 ;
      RECT 917.420 1.400 917.700 980.000 ;
      RECT 919.660 1.400 919.940 980.000 ;
      RECT 921.900 1.400 922.180 980.000 ;
      RECT 924.140 1.400 924.420 980.000 ;
      RECT 926.380 1.400 926.660 980.000 ;
      RECT 928.620 1.400 928.900 980.000 ;
      RECT 930.860 1.400 931.140 980.000 ;
      RECT 933.100 1.400 933.380 980.000 ;
      RECT 935.340 1.400 935.620 980.000 ;
      RECT 937.580 1.400 937.860 980.000 ;
      RECT 939.820 1.400 940.100 980.000 ;
      RECT 942.060 1.400 942.340 980.000 ;
      RECT 944.300 1.400 944.580 980.000 ;
      RECT 946.540 1.400 946.820 980.000 ;
      RECT 948.780 1.400 949.060 980.000 ;
      RECT 951.020 1.400 951.300 980.000 ;
      RECT 953.260 1.400 953.540 980.000 ;
      RECT 955.500 1.400 955.780 980.000 ;
      RECT 957.740 1.400 958.020 980.000 ;
      RECT 959.980 1.400 960.260 980.000 ;
      RECT 962.220 1.400 962.500 980.000 ;
      RECT 964.460 1.400 964.740 980.000 ;
      RECT 966.700 1.400 966.980 980.000 ;
      RECT 968.940 1.400 969.220 980.000 ;
      RECT 971.180 1.400 971.460 980.000 ;
      RECT 973.420 1.400 973.700 980.000 ;
      RECT 975.660 1.400 975.940 980.000 ;
      RECT 977.900 1.400 978.180 980.000 ;
      RECT 980.140 1.400 980.420 980.000 ;
      RECT 982.380 1.400 982.660 980.000 ;
      RECT 984.620 1.400 984.900 980.000 ;
      RECT 986.860 1.400 987.140 980.000 ;
      RECT 989.100 1.400 989.380 980.000 ;
      RECT 991.340 1.400 991.620 980.000 ;
      RECT 993.580 1.400 993.860 980.000 ;
      RECT 995.820 1.400 996.100 980.000 ;
      RECT 998.060 1.400 998.340 980.000 ;
      RECT 1000.300 1.400 1000.580 980.000 ;
      RECT 1002.540 1.400 1002.820 980.000 ;
      RECT 1004.780 1.400 1005.060 980.000 ;
      RECT 1007.020 1.400 1007.300 980.000 ;
      RECT 1009.260 1.400 1009.540 980.000 ;
      RECT 1011.500 1.400 1011.780 980.000 ;
      RECT 1013.740 1.400 1014.020 980.000 ;
      RECT 1015.980 1.400 1016.260 980.000 ;
      RECT 1018.220 1.400 1018.500 980.000 ;
      RECT 1020.460 1.400 1020.740 980.000 ;
      RECT 1022.700 1.400 1022.980 980.000 ;
      RECT 1024.940 1.400 1025.220 980.000 ;
      RECT 1027.180 1.400 1027.460 980.000 ;
      RECT 1029.420 1.400 1029.700 980.000 ;
      RECT 1031.660 1.400 1031.940 980.000 ;
      RECT 1033.900 1.400 1034.180 980.000 ;
      RECT 1036.140 1.400 1036.420 980.000 ;
      RECT 1038.380 1.400 1038.660 980.000 ;
      RECT 1040.620 1.400 1040.900 980.000 ;
      RECT 1042.860 1.400 1043.140 980.000 ;
      RECT 1045.100 1.400 1045.380 980.000 ;
      RECT 1047.340 1.400 1047.620 980.000 ;
      RECT 1049.580 1.400 1049.860 980.000 ;
      RECT 1051.820 1.400 1052.100 980.000 ;
      RECT 1054.060 1.400 1054.340 980.000 ;
      RECT 1056.300 1.400 1056.580 980.000 ;
      RECT 1058.540 1.400 1058.820 980.000 ;
      RECT 1060.780 1.400 1061.060 980.000 ;
      RECT 1063.020 1.400 1063.300 980.000 ;
      RECT 1065.260 1.400 1065.540 980.000 ;
      RECT 1067.500 1.400 1067.780 980.000 ;
      RECT 1069.740 1.400 1070.020 980.000 ;
      RECT 1071.980 1.400 1072.260 980.000 ;
      RECT 1074.220 1.400 1074.500 980.000 ;
      RECT 1076.460 1.400 1076.740 980.000 ;
      RECT 1078.700 1.400 1078.980 980.000 ;
      RECT 1080.940 1.400 1081.220 980.000 ;
      RECT 1083.180 1.400 1083.460 980.000 ;
      RECT 1085.420 1.400 1085.700 980.000 ;
      RECT 1087.660 1.400 1087.940 980.000 ;
      RECT 1089.900 1.400 1090.180 980.000 ;
      RECT 1092.140 1.400 1092.420 980.000 ;
      RECT 1094.380 1.400 1094.660 980.000 ;
      RECT 1096.620 1.400 1096.900 980.000 ;
      RECT 1098.860 1.400 1099.140 980.000 ;
      RECT 1101.100 1.400 1101.380 980.000 ;
      RECT 1103.340 1.400 1103.620 980.000 ;
      RECT 1105.580 1.400 1105.860 980.000 ;
      RECT 1107.820 1.400 1108.100 980.000 ;
      RECT 1110.060 1.400 1110.340 980.000 ;
      RECT 1112.300 1.400 1112.580 980.000 ;
      RECT 1114.540 1.400 1114.820 980.000 ;
      RECT 1116.780 1.400 1117.060 980.000 ;
      RECT 1119.020 1.400 1119.300 980.000 ;
      RECT 1121.260 1.400 1121.540 980.000 ;
      RECT 1123.500 1.400 1123.780 980.000 ;
      RECT 1125.740 1.400 1126.020 980.000 ;
      RECT 1127.980 1.400 1128.260 980.000 ;
      RECT 1130.220 1.400 1130.500 980.000 ;
      RECT 1132.460 1.400 1132.740 980.000 ;
      RECT 1134.700 1.400 1134.980 980.000 ;
      RECT 1136.940 1.400 1137.220 980.000 ;
      RECT 1139.180 1.400 1139.460 980.000 ;
      RECT 1141.420 1.400 1141.700 980.000 ;
      RECT 1143.660 1.400 1143.940 980.000 ;
      RECT 1145.900 1.400 1146.180 980.000 ;
      RECT 1148.140 1.400 1148.420 980.000 ;
      RECT 1150.380 1.400 1150.660 980.000 ;
      RECT 1152.620 1.400 1152.900 980.000 ;
      RECT 1154.860 1.400 1155.140 980.000 ;
      RECT 1157.100 1.400 1157.380 980.000 ;
      RECT 1159.340 1.400 1159.620 980.000 ;
      RECT 1161.580 1.400 1161.860 980.000 ;
      RECT 1163.820 1.400 1164.100 980.000 ;
      RECT 1166.060 1.400 1166.340 980.000 ;
      RECT 1168.300 1.400 1168.580 980.000 ;
      RECT 1170.540 1.400 1170.820 980.000 ;
      RECT 1172.780 1.400 1173.060 980.000 ;
      RECT 1175.020 1.400 1175.300 980.000 ;
      RECT 1177.260 1.400 1177.540 980.000 ;
      RECT 1179.500 1.400 1179.780 980.000 ;
      RECT 1181.740 1.400 1182.020 980.000 ;
      RECT 1183.980 1.400 1184.260 980.000 ;
      RECT 1186.220 1.400 1186.500 980.000 ;
      RECT 1188.460 1.400 1188.740 980.000 ;
      RECT 1190.700 1.400 1190.980 980.000 ;
      RECT 1192.940 1.400 1193.220 980.000 ;
      RECT 1195.180 1.400 1195.460 980.000 ;
      RECT 1197.420 1.400 1197.700 980.000 ;
      RECT 1199.660 1.400 1199.940 980.000 ;
      RECT 1201.900 1.400 1202.180 980.000 ;
      RECT 1204.140 1.400 1204.420 980.000 ;
      RECT 1206.380 1.400 1206.660 980.000 ;
      RECT 1208.620 1.400 1208.900 980.000 ;
      RECT 1210.860 1.400 1211.140 980.000 ;
      RECT 1213.100 1.400 1213.380 980.000 ;
      RECT 1215.340 1.400 1215.620 980.000 ;
      RECT 1217.580 1.400 1217.860 980.000 ;
      RECT 1219.820 1.400 1220.100 980.000 ;
      RECT 1222.060 1.400 1222.340 980.000 ;
      RECT 1224.300 1.400 1224.580 980.000 ;
      RECT 1226.540 1.400 1226.820 980.000 ;
      RECT 1228.780 1.400 1229.060 980.000 ;
      RECT 1231.020 1.400 1231.300 980.000 ;
      RECT 1233.260 1.400 1233.540 980.000 ;
      RECT 1235.500 1.400 1235.780 980.000 ;
      RECT 1237.740 1.400 1238.020 980.000 ;
      RECT 1239.980 1.400 1240.260 980.000 ;
      RECT 1242.220 1.400 1242.500 980.000 ;
      RECT 1244.460 1.400 1244.740 980.000 ;
      RECT 1246.700 1.400 1246.980 980.000 ;
      RECT 1248.940 1.400 1249.220 980.000 ;
      RECT 1251.180 1.400 1251.460 980.000 ;
      RECT 1253.420 1.400 1253.700 980.000 ;
      RECT 1255.660 1.400 1255.940 980.000 ;
      RECT 1257.900 1.400 1258.180 980.000 ;
      RECT 1260.140 1.400 1260.420 980.000 ;
      RECT 1262.380 1.400 1262.660 980.000 ;
      RECT 1264.620 1.400 1264.900 980.000 ;
      RECT 1266.860 1.400 1267.140 980.000 ;
      RECT 1269.100 1.400 1269.380 980.000 ;
      RECT 1271.340 1.400 1271.620 980.000 ;
      RECT 1273.580 1.400 1273.860 980.000 ;
      RECT 1275.820 1.400 1276.100 980.000 ;
      RECT 1278.060 1.400 1278.340 980.000 ;
      RECT 1280.300 1.400 1280.580 980.000 ;
      RECT 1282.540 1.400 1282.820 980.000 ;
      RECT 1284.780 1.400 1285.060 980.000 ;
      RECT 1287.020 1.400 1287.300 980.000 ;
      RECT 1289.260 1.400 1289.540 980.000 ;
      RECT 1291.500 1.400 1291.780 980.000 ;
      RECT 1293.740 1.400 1294.020 980.000 ;
      RECT 1295.980 1.400 1296.260 980.000 ;
      RECT 1298.220 1.400 1298.500 980.000 ;
      RECT 1300.460 1.400 1300.740 980.000 ;
      RECT 1302.700 1.400 1302.980 980.000 ;
      RECT 1304.940 1.400 1305.220 980.000 ;
      RECT 1307.180 1.400 1307.460 980.000 ;
      RECT 1309.420 1.400 1309.700 980.000 ;
      RECT 1311.660 1.400 1311.940 980.000 ;
      RECT 1313.900 1.400 1314.180 980.000 ;
      RECT 1316.140 1.400 1316.420 980.000 ;
      RECT 1318.380 1.400 1318.660 980.000 ;
      RECT 1320.620 1.400 1320.900 980.000 ;
      RECT 1322.860 1.400 1323.140 980.000 ;
      RECT 1325.100 1.400 1325.380 980.000 ;
      RECT 1327.340 1.400 1327.620 980.000 ;
      RECT 1329.580 1.400 1329.860 980.000 ;
      RECT 1331.820 1.400 1332.100 980.000 ;
      RECT 1334.060 1.400 1334.340 980.000 ;
      RECT 1336.300 1.400 1336.580 980.000 ;
      RECT 1338.540 1.400 1338.820 980.000 ;
      RECT 1340.780 1.400 1341.060 980.000 ;
      RECT 1343.020 1.400 1343.300 980.000 ;
      RECT 1345.260 1.400 1345.540 980.000 ;
      RECT 1347.500 1.400 1347.780 980.000 ;
      RECT 1349.740 1.400 1350.020 980.000 ;
      RECT 1351.980 1.400 1352.260 980.000 ;
      RECT 1354.220 1.400 1354.500 980.000 ;
      RECT 1356.460 1.400 1356.740 980.000 ;
      RECT 1358.700 1.400 1358.980 980.000 ;
      RECT 1360.940 1.400 1361.220 980.000 ;
      RECT 1363.180 1.400 1363.460 980.000 ;
      RECT 1365.420 1.400 1365.700 980.000 ;
      RECT 1367.660 1.400 1367.940 980.000 ;
      RECT 1369.900 1.400 1370.180 980.000 ;
      RECT 1372.140 1.400 1372.420 980.000 ;
      RECT 1374.380 1.400 1374.660 980.000 ;
      RECT 1376.620 1.400 1376.900 980.000 ;
      RECT 1378.860 1.400 1379.140 980.000 ;
      RECT 1381.100 1.400 1381.380 980.000 ;
      RECT 1383.340 1.400 1383.620 980.000 ;
      RECT 1385.580 1.400 1385.860 980.000 ;
      RECT 1387.820 1.400 1388.100 980.000 ;
      RECT 1390.060 1.400 1390.340 980.000 ;
      RECT 1392.300 1.400 1392.580 980.000 ;
      RECT 1394.540 1.400 1394.820 980.000 ;
      RECT 1396.780 1.400 1397.060 980.000 ;
      RECT 1399.020 1.400 1399.300 980.000 ;
      RECT 1401.260 1.400 1401.540 980.000 ;
      RECT 1403.500 1.400 1403.780 980.000 ;
      RECT 1405.740 1.400 1406.020 980.000 ;
      RECT 1407.980 1.400 1408.260 980.000 ;
      RECT 1410.220 1.400 1410.500 980.000 ;
      RECT 1412.460 1.400 1412.740 980.000 ;
      RECT 1414.700 1.400 1414.980 980.000 ;
      RECT 1416.940 1.400 1417.220 980.000 ;
      RECT 1419.180 1.400 1419.460 980.000 ;
      RECT 1421.420 1.400 1421.700 980.000 ;
      RECT 1423.660 1.400 1423.940 980.000 ;
      RECT 1425.900 1.400 1426.180 980.000 ;
      RECT 1428.140 1.400 1428.420 980.000 ;
      RECT 1430.380 1.400 1430.660 980.000 ;
      RECT 1432.620 1.400 1432.900 980.000 ;
      RECT 1434.860 1.400 1435.140 980.000 ;
      RECT 1437.100 1.400 1437.380 980.000 ;
      RECT 1439.340 1.400 1439.620 980.000 ;
      RECT 1441.580 1.400 1441.860 980.000 ;
      RECT 1443.820 1.400 1444.100 980.000 ;
      RECT 1446.060 1.400 1446.340 980.000 ;
      RECT 1448.300 1.400 1448.580 980.000 ;
      RECT 1450.540 1.400 1450.820 980.000 ;
      RECT 1452.780 1.400 1453.060 980.000 ;
      RECT 1455.020 1.400 1455.300 980.000 ;
      RECT 1457.260 1.400 1457.540 980.000 ;
      RECT 1459.500 1.400 1459.780 980.000 ;
      RECT 1461.740 1.400 1462.020 980.000 ;
      RECT 1463.980 1.400 1464.260 980.000 ;
      RECT 1466.220 1.400 1466.500 980.000 ;
      RECT 1468.460 1.400 1468.740 980.000 ;
      RECT 1470.700 1.400 1470.980 980.000 ;
      RECT 1472.940 1.400 1473.220 980.000 ;
      RECT 1475.180 1.400 1475.460 980.000 ;
      RECT 1477.420 1.400 1477.700 980.000 ;
      RECT 1479.660 1.400 1479.940 980.000 ;
      RECT 1481.900 1.400 1482.180 980.000 ;
      RECT 1484.140 1.400 1484.420 980.000 ;
      RECT 1486.380 1.400 1486.660 980.000 ;
      RECT 1488.620 1.400 1488.900 980.000 ;
      RECT 1490.860 1.400 1491.140 980.000 ;
      RECT 1493.100 1.400 1493.380 980.000 ;
      RECT 1495.340 1.400 1495.620 980.000 ;
      RECT 1497.580 1.400 1497.860 980.000 ;
      RECT 1499.820 1.400 1500.100 980.000 ;
      RECT 1502.060 1.400 1502.340 980.000 ;
      RECT 1504.300 1.400 1504.580 980.000 ;
      RECT 1506.540 1.400 1506.820 980.000 ;
      RECT 1508.780 1.400 1509.060 980.000 ;
      RECT 1511.020 1.400 1511.300 980.000 ;
      RECT 1513.260 1.400 1513.540 980.000 ;
      RECT 1515.500 1.400 1515.780 980.000 ;
      RECT 1517.740 1.400 1518.020 980.000 ;
      RECT 1519.980 1.400 1520.260 980.000 ;
      RECT 1522.220 1.400 1522.500 980.000 ;
      RECT 1524.460 1.400 1524.740 980.000 ;
      RECT 1526.700 1.400 1526.980 980.000 ;
      RECT 1528.940 1.400 1529.220 980.000 ;
      RECT 1531.180 1.400 1531.460 980.000 ;
      RECT 1533.420 1.400 1533.700 980.000 ;
      RECT 1535.660 1.400 1535.940 980.000 ;
      RECT 1537.900 1.400 1538.180 980.000 ;
      RECT 1540.140 1.400 1540.420 980.000 ;
      RECT 1542.380 1.400 1542.660 980.000 ;
      RECT 1544.620 1.400 1544.900 980.000 ;
      RECT 1546.860 1.400 1547.140 980.000 ;
      RECT 1549.100 1.400 1549.380 980.000 ;
      RECT 1551.340 1.400 1551.620 980.000 ;
      RECT 1553.580 1.400 1553.860 980.000 ;
      RECT 1555.820 1.400 1556.100 980.000 ;
      RECT 1558.060 1.400 1558.340 980.000 ;
      RECT 1560.300 1.400 1560.580 980.000 ;
      RECT 1562.540 1.400 1562.820 980.000 ;
      RECT 1564.780 1.400 1565.060 980.000 ;
      RECT 1567.020 1.400 1567.300 980.000 ;
      RECT 1569.260 1.400 1569.540 980.000 ;
      RECT 1571.500 1.400 1571.780 980.000 ;
      RECT 1573.740 1.400 1574.020 980.000 ;
      RECT 1575.980 1.400 1576.260 980.000 ;
      RECT 1578.220 1.400 1578.500 980.000 ;
      RECT 1580.460 1.400 1580.740 980.000 ;
      RECT 1582.700 1.400 1582.980 980.000 ;
      RECT 1584.940 1.400 1585.220 980.000 ;
      RECT 1587.180 1.400 1587.460 980.000 ;
      RECT 1589.420 1.400 1589.700 980.000 ;
      RECT 1591.660 1.400 1591.940 980.000 ;
      RECT 1593.900 1.400 1594.180 980.000 ;
      RECT 1596.140 1.400 1596.420 980.000 ;
      RECT 1598.380 1.400 1598.660 980.000 ;
      RECT 1600.620 1.400 1600.900 980.000 ;
      RECT 1602.860 1.400 1603.140 980.000 ;
      RECT 1605.100 1.400 1605.380 980.000 ;
      RECT 1607.340 1.400 1607.620 980.000 ;
      RECT 1609.580 1.400 1609.860 980.000 ;
      RECT 1611.820 1.400 1612.100 980.000 ;
      RECT 1614.060 1.400 1614.340 980.000 ;
      RECT 1616.300 1.400 1616.580 980.000 ;
      RECT 1618.540 1.400 1618.820 980.000 ;
      RECT 1620.780 1.400 1621.060 980.000 ;
      RECT 1623.020 1.400 1623.300 980.000 ;
      RECT 1625.260 1.400 1625.540 980.000 ;
      RECT 1627.500 1.400 1627.780 980.000 ;
      RECT 1629.740 1.400 1630.020 980.000 ;
      RECT 1631.980 1.400 1632.260 980.000 ;
      RECT 1634.220 1.400 1634.500 980.000 ;
      RECT 1636.460 1.400 1636.740 980.000 ;
      RECT 1638.700 1.400 1638.980 980.000 ;
      RECT 1640.940 1.400 1641.220 980.000 ;
      RECT 1643.180 1.400 1643.460 980.000 ;
      RECT 1645.420 1.400 1645.700 980.000 ;
      RECT 1647.660 1.400 1647.940 980.000 ;
      RECT 1649.900 1.400 1650.180 980.000 ;
      RECT 1652.140 1.400 1652.420 980.000 ;
      RECT 1654.380 1.400 1654.660 980.000 ;
      RECT 1656.620 1.400 1656.900 980.000 ;
      RECT 1658.860 1.400 1659.140 980.000 ;
      RECT 1661.100 1.400 1661.380 980.000 ;
      RECT 1663.340 1.400 1663.620 980.000 ;
      RECT 1665.580 1.400 1665.860 980.000 ;
      RECT 1667.820 1.400 1668.100 980.000 ;
      RECT 1670.060 1.400 1670.340 980.000 ;
      RECT 1672.300 1.400 1672.580 980.000 ;
      RECT 1674.540 1.400 1674.820 980.000 ;
      RECT 1676.780 1.400 1677.060 980.000 ;
      RECT 1679.020 1.400 1679.300 980.000 ;
      RECT 1681.260 1.400 1681.540 980.000 ;
      RECT 1683.500 1.400 1683.780 980.000 ;
      RECT 1685.740 1.400 1686.020 980.000 ;
      RECT 1687.980 1.400 1688.260 980.000 ;
      RECT 1690.220 1.400 1690.500 980.000 ;
      RECT 1692.460 1.400 1692.740 980.000 ;
      RECT 1694.700 1.400 1694.980 980.000 ;
      RECT 1696.940 1.400 1697.220 980.000 ;
      RECT 1699.180 1.400 1699.460 980.000 ;
      RECT 1701.420 1.400 1701.700 980.000 ;
      RECT 1703.660 1.400 1703.940 980.000 ;
      RECT 1705.900 1.400 1706.180 980.000 ;
      RECT 1708.140 1.400 1708.420 980.000 ;
      RECT 1710.380 1.400 1710.660 980.000 ;
      RECT 1712.620 1.400 1712.900 980.000 ;
      RECT 1714.860 1.400 1715.140 980.000 ;
      RECT 1717.100 1.400 1717.380 980.000 ;
      RECT 1719.340 1.400 1719.620 980.000 ;
      RECT 1721.580 1.400 1721.860 980.000 ;
      RECT 1723.820 1.400 1724.100 980.000 ;
      RECT 1726.060 1.400 1726.340 980.000 ;
      RECT 1728.300 1.400 1728.580 980.000 ;
      RECT 1730.540 1.400 1730.820 980.000 ;
      RECT 1732.780 1.400 1733.060 980.000 ;
      RECT 1735.020 1.400 1735.300 980.000 ;
      RECT 1737.260 1.400 1737.540 980.000 ;
      RECT 1739.500 1.400 1739.780 980.000 ;
      RECT 1741.740 1.400 1742.020 980.000 ;
      RECT 1743.980 1.400 1744.260 980.000 ;
      RECT 1746.220 1.400 1746.500 980.000 ;
      RECT 1748.460 1.400 1748.740 980.000 ;
      RECT 1750.700 1.400 1750.980 980.000 ;
      RECT 1752.940 1.400 1753.220 980.000 ;
      RECT 1755.180 1.400 1755.460 980.000 ;
      RECT 1757.420 1.400 1757.700 980.000 ;
      RECT 1759.660 1.400 1759.940 980.000 ;
      RECT 1761.900 1.400 1762.180 980.000 ;
      RECT 1764.140 1.400 1764.420 980.000 ;
      RECT 1766.380 1.400 1766.660 980.000 ;
      RECT 1768.620 1.400 1768.900 980.000 ;
      RECT 1770.860 1.400 1771.140 980.000 ;
      RECT 1773.100 1.400 1773.380 980.000 ;
      RECT 1775.340 1.400 1775.620 980.000 ;
      RECT 1777.580 1.400 1777.860 980.000 ;
      RECT 1779.820 1.400 1780.100 980.000 ;
      RECT 1782.060 1.400 1782.340 980.000 ;
      RECT 1784.300 1.400 1784.580 980.000 ;
      RECT 1786.540 1.400 1786.820 980.000 ;
      RECT 1788.780 1.400 1789.060 980.000 ;
      RECT 1791.020 1.400 1791.300 980.000 ;
      RECT 1793.260 1.400 1793.540 980.000 ;
      RECT 1795.500 1.400 1795.780 980.000 ;
      RECT 1797.740 1.400 1798.020 980.000 ;
      RECT 1799.980 1.400 1800.260 980.000 ;
      RECT 1802.220 1.400 1802.500 980.000 ;
      RECT 1804.460 1.400 1804.740 980.000 ;
      RECT 1806.700 1.400 1806.980 980.000 ;
      RECT 1808.940 1.400 1809.220 980.000 ;
      RECT 1811.180 1.400 1811.460 980.000 ;
      RECT 1813.420 1.400 1813.700 980.000 ;
      RECT 1815.660 1.400 1815.940 980.000 ;
      RECT 1817.900 1.400 1818.180 980.000 ;
      RECT 1820.140 1.400 1820.420 980.000 ;
      RECT 1822.380 1.400 1822.660 980.000 ;
      RECT 1824.620 1.400 1824.900 980.000 ;
      RECT 1826.860 1.400 1827.140 980.000 ;
      RECT 1829.100 1.400 1829.380 980.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 980.000 ;
      RECT 4.620 1.400 4.900 980.000 ;
      RECT 6.860 1.400 7.140 980.000 ;
      RECT 9.100 1.400 9.380 980.000 ;
      RECT 11.340 1.400 11.620 980.000 ;
      RECT 13.580 1.400 13.860 980.000 ;
      RECT 15.820 1.400 16.100 980.000 ;
      RECT 18.060 1.400 18.340 980.000 ;
      RECT 20.300 1.400 20.580 980.000 ;
      RECT 22.540 1.400 22.820 980.000 ;
      RECT 24.780 1.400 25.060 980.000 ;
      RECT 27.020 1.400 27.300 980.000 ;
      RECT 29.260 1.400 29.540 980.000 ;
      RECT 31.500 1.400 31.780 980.000 ;
      RECT 33.740 1.400 34.020 980.000 ;
      RECT 35.980 1.400 36.260 980.000 ;
      RECT 38.220 1.400 38.500 980.000 ;
      RECT 40.460 1.400 40.740 980.000 ;
      RECT 42.700 1.400 42.980 980.000 ;
      RECT 44.940 1.400 45.220 980.000 ;
      RECT 47.180 1.400 47.460 980.000 ;
      RECT 49.420 1.400 49.700 980.000 ;
      RECT 51.660 1.400 51.940 980.000 ;
      RECT 53.900 1.400 54.180 980.000 ;
      RECT 56.140 1.400 56.420 980.000 ;
      RECT 58.380 1.400 58.660 980.000 ;
      RECT 60.620 1.400 60.900 980.000 ;
      RECT 62.860 1.400 63.140 980.000 ;
      RECT 65.100 1.400 65.380 980.000 ;
      RECT 67.340 1.400 67.620 980.000 ;
      RECT 69.580 1.400 69.860 980.000 ;
      RECT 71.820 1.400 72.100 980.000 ;
      RECT 74.060 1.400 74.340 980.000 ;
      RECT 76.300 1.400 76.580 980.000 ;
      RECT 78.540 1.400 78.820 980.000 ;
      RECT 80.780 1.400 81.060 980.000 ;
      RECT 83.020 1.400 83.300 980.000 ;
      RECT 85.260 1.400 85.540 980.000 ;
      RECT 87.500 1.400 87.780 980.000 ;
      RECT 89.740 1.400 90.020 980.000 ;
      RECT 91.980 1.400 92.260 980.000 ;
      RECT 94.220 1.400 94.500 980.000 ;
      RECT 96.460 1.400 96.740 980.000 ;
      RECT 98.700 1.400 98.980 980.000 ;
      RECT 100.940 1.400 101.220 980.000 ;
      RECT 103.180 1.400 103.460 980.000 ;
      RECT 105.420 1.400 105.700 980.000 ;
      RECT 107.660 1.400 107.940 980.000 ;
      RECT 109.900 1.400 110.180 980.000 ;
      RECT 112.140 1.400 112.420 980.000 ;
      RECT 114.380 1.400 114.660 980.000 ;
      RECT 116.620 1.400 116.900 980.000 ;
      RECT 118.860 1.400 119.140 980.000 ;
      RECT 121.100 1.400 121.380 980.000 ;
      RECT 123.340 1.400 123.620 980.000 ;
      RECT 125.580 1.400 125.860 980.000 ;
      RECT 127.820 1.400 128.100 980.000 ;
      RECT 130.060 1.400 130.340 980.000 ;
      RECT 132.300 1.400 132.580 980.000 ;
      RECT 134.540 1.400 134.820 980.000 ;
      RECT 136.780 1.400 137.060 980.000 ;
      RECT 139.020 1.400 139.300 980.000 ;
      RECT 141.260 1.400 141.540 980.000 ;
      RECT 143.500 1.400 143.780 980.000 ;
      RECT 145.740 1.400 146.020 980.000 ;
      RECT 147.980 1.400 148.260 980.000 ;
      RECT 150.220 1.400 150.500 980.000 ;
      RECT 152.460 1.400 152.740 980.000 ;
      RECT 154.700 1.400 154.980 980.000 ;
      RECT 156.940 1.400 157.220 980.000 ;
      RECT 159.180 1.400 159.460 980.000 ;
      RECT 161.420 1.400 161.700 980.000 ;
      RECT 163.660 1.400 163.940 980.000 ;
      RECT 165.900 1.400 166.180 980.000 ;
      RECT 168.140 1.400 168.420 980.000 ;
      RECT 170.380 1.400 170.660 980.000 ;
      RECT 172.620 1.400 172.900 980.000 ;
      RECT 174.860 1.400 175.140 980.000 ;
      RECT 177.100 1.400 177.380 980.000 ;
      RECT 179.340 1.400 179.620 980.000 ;
      RECT 181.580 1.400 181.860 980.000 ;
      RECT 183.820 1.400 184.100 980.000 ;
      RECT 186.060 1.400 186.340 980.000 ;
      RECT 188.300 1.400 188.580 980.000 ;
      RECT 190.540 1.400 190.820 980.000 ;
      RECT 192.780 1.400 193.060 980.000 ;
      RECT 195.020 1.400 195.300 980.000 ;
      RECT 197.260 1.400 197.540 980.000 ;
      RECT 199.500 1.400 199.780 980.000 ;
      RECT 201.740 1.400 202.020 980.000 ;
      RECT 203.980 1.400 204.260 980.000 ;
      RECT 206.220 1.400 206.500 980.000 ;
      RECT 208.460 1.400 208.740 980.000 ;
      RECT 210.700 1.400 210.980 980.000 ;
      RECT 212.940 1.400 213.220 980.000 ;
      RECT 215.180 1.400 215.460 980.000 ;
      RECT 217.420 1.400 217.700 980.000 ;
      RECT 219.660 1.400 219.940 980.000 ;
      RECT 221.900 1.400 222.180 980.000 ;
      RECT 224.140 1.400 224.420 980.000 ;
      RECT 226.380 1.400 226.660 980.000 ;
      RECT 228.620 1.400 228.900 980.000 ;
      RECT 230.860 1.400 231.140 980.000 ;
      RECT 233.100 1.400 233.380 980.000 ;
      RECT 235.340 1.400 235.620 980.000 ;
      RECT 237.580 1.400 237.860 980.000 ;
      RECT 239.820 1.400 240.100 980.000 ;
      RECT 242.060 1.400 242.340 980.000 ;
      RECT 244.300 1.400 244.580 980.000 ;
      RECT 246.540 1.400 246.820 980.000 ;
      RECT 248.780 1.400 249.060 980.000 ;
      RECT 251.020 1.400 251.300 980.000 ;
      RECT 253.260 1.400 253.540 980.000 ;
      RECT 255.500 1.400 255.780 980.000 ;
      RECT 257.740 1.400 258.020 980.000 ;
      RECT 259.980 1.400 260.260 980.000 ;
      RECT 262.220 1.400 262.500 980.000 ;
      RECT 264.460 1.400 264.740 980.000 ;
      RECT 266.700 1.400 266.980 980.000 ;
      RECT 268.940 1.400 269.220 980.000 ;
      RECT 271.180 1.400 271.460 980.000 ;
      RECT 273.420 1.400 273.700 980.000 ;
      RECT 275.660 1.400 275.940 980.000 ;
      RECT 277.900 1.400 278.180 980.000 ;
      RECT 280.140 1.400 280.420 980.000 ;
      RECT 282.380 1.400 282.660 980.000 ;
      RECT 284.620 1.400 284.900 980.000 ;
      RECT 286.860 1.400 287.140 980.000 ;
      RECT 289.100 1.400 289.380 980.000 ;
      RECT 291.340 1.400 291.620 980.000 ;
      RECT 293.580 1.400 293.860 980.000 ;
      RECT 295.820 1.400 296.100 980.000 ;
      RECT 298.060 1.400 298.340 980.000 ;
      RECT 300.300 1.400 300.580 980.000 ;
      RECT 302.540 1.400 302.820 980.000 ;
      RECT 304.780 1.400 305.060 980.000 ;
      RECT 307.020 1.400 307.300 980.000 ;
      RECT 309.260 1.400 309.540 980.000 ;
      RECT 311.500 1.400 311.780 980.000 ;
      RECT 313.740 1.400 314.020 980.000 ;
      RECT 315.980 1.400 316.260 980.000 ;
      RECT 318.220 1.400 318.500 980.000 ;
      RECT 320.460 1.400 320.740 980.000 ;
      RECT 322.700 1.400 322.980 980.000 ;
      RECT 324.940 1.400 325.220 980.000 ;
      RECT 327.180 1.400 327.460 980.000 ;
      RECT 329.420 1.400 329.700 980.000 ;
      RECT 331.660 1.400 331.940 980.000 ;
      RECT 333.900 1.400 334.180 980.000 ;
      RECT 336.140 1.400 336.420 980.000 ;
      RECT 338.380 1.400 338.660 980.000 ;
      RECT 340.620 1.400 340.900 980.000 ;
      RECT 342.860 1.400 343.140 980.000 ;
      RECT 345.100 1.400 345.380 980.000 ;
      RECT 347.340 1.400 347.620 980.000 ;
      RECT 349.580 1.400 349.860 980.000 ;
      RECT 351.820 1.400 352.100 980.000 ;
      RECT 354.060 1.400 354.340 980.000 ;
      RECT 356.300 1.400 356.580 980.000 ;
      RECT 358.540 1.400 358.820 980.000 ;
      RECT 360.780 1.400 361.060 980.000 ;
      RECT 363.020 1.400 363.300 980.000 ;
      RECT 365.260 1.400 365.540 980.000 ;
      RECT 367.500 1.400 367.780 980.000 ;
      RECT 369.740 1.400 370.020 980.000 ;
      RECT 371.980 1.400 372.260 980.000 ;
      RECT 374.220 1.400 374.500 980.000 ;
      RECT 376.460 1.400 376.740 980.000 ;
      RECT 378.700 1.400 378.980 980.000 ;
      RECT 380.940 1.400 381.220 980.000 ;
      RECT 383.180 1.400 383.460 980.000 ;
      RECT 385.420 1.400 385.700 980.000 ;
      RECT 387.660 1.400 387.940 980.000 ;
      RECT 389.900 1.400 390.180 980.000 ;
      RECT 392.140 1.400 392.420 980.000 ;
      RECT 394.380 1.400 394.660 980.000 ;
      RECT 396.620 1.400 396.900 980.000 ;
      RECT 398.860 1.400 399.140 980.000 ;
      RECT 401.100 1.400 401.380 980.000 ;
      RECT 403.340 1.400 403.620 980.000 ;
      RECT 405.580 1.400 405.860 980.000 ;
      RECT 407.820 1.400 408.100 980.000 ;
      RECT 410.060 1.400 410.340 980.000 ;
      RECT 412.300 1.400 412.580 980.000 ;
      RECT 414.540 1.400 414.820 980.000 ;
      RECT 416.780 1.400 417.060 980.000 ;
      RECT 419.020 1.400 419.300 980.000 ;
      RECT 421.260 1.400 421.540 980.000 ;
      RECT 423.500 1.400 423.780 980.000 ;
      RECT 425.740 1.400 426.020 980.000 ;
      RECT 427.980 1.400 428.260 980.000 ;
      RECT 430.220 1.400 430.500 980.000 ;
      RECT 432.460 1.400 432.740 980.000 ;
      RECT 434.700 1.400 434.980 980.000 ;
      RECT 436.940 1.400 437.220 980.000 ;
      RECT 439.180 1.400 439.460 980.000 ;
      RECT 441.420 1.400 441.700 980.000 ;
      RECT 443.660 1.400 443.940 980.000 ;
      RECT 445.900 1.400 446.180 980.000 ;
      RECT 448.140 1.400 448.420 980.000 ;
      RECT 450.380 1.400 450.660 980.000 ;
      RECT 452.620 1.400 452.900 980.000 ;
      RECT 454.860 1.400 455.140 980.000 ;
      RECT 457.100 1.400 457.380 980.000 ;
      RECT 459.340 1.400 459.620 980.000 ;
      RECT 461.580 1.400 461.860 980.000 ;
      RECT 463.820 1.400 464.100 980.000 ;
      RECT 466.060 1.400 466.340 980.000 ;
      RECT 468.300 1.400 468.580 980.000 ;
      RECT 470.540 1.400 470.820 980.000 ;
      RECT 472.780 1.400 473.060 980.000 ;
      RECT 475.020 1.400 475.300 980.000 ;
      RECT 477.260 1.400 477.540 980.000 ;
      RECT 479.500 1.400 479.780 980.000 ;
      RECT 481.740 1.400 482.020 980.000 ;
      RECT 483.980 1.400 484.260 980.000 ;
      RECT 486.220 1.400 486.500 980.000 ;
      RECT 488.460 1.400 488.740 980.000 ;
      RECT 490.700 1.400 490.980 980.000 ;
      RECT 492.940 1.400 493.220 980.000 ;
      RECT 495.180 1.400 495.460 980.000 ;
      RECT 497.420 1.400 497.700 980.000 ;
      RECT 499.660 1.400 499.940 980.000 ;
      RECT 501.900 1.400 502.180 980.000 ;
      RECT 504.140 1.400 504.420 980.000 ;
      RECT 506.380 1.400 506.660 980.000 ;
      RECT 508.620 1.400 508.900 980.000 ;
      RECT 510.860 1.400 511.140 980.000 ;
      RECT 513.100 1.400 513.380 980.000 ;
      RECT 515.340 1.400 515.620 980.000 ;
      RECT 517.580 1.400 517.860 980.000 ;
      RECT 519.820 1.400 520.100 980.000 ;
      RECT 522.060 1.400 522.340 980.000 ;
      RECT 524.300 1.400 524.580 980.000 ;
      RECT 526.540 1.400 526.820 980.000 ;
      RECT 528.780 1.400 529.060 980.000 ;
      RECT 531.020 1.400 531.300 980.000 ;
      RECT 533.260 1.400 533.540 980.000 ;
      RECT 535.500 1.400 535.780 980.000 ;
      RECT 537.740 1.400 538.020 980.000 ;
      RECT 539.980 1.400 540.260 980.000 ;
      RECT 542.220 1.400 542.500 980.000 ;
      RECT 544.460 1.400 544.740 980.000 ;
      RECT 546.700 1.400 546.980 980.000 ;
      RECT 548.940 1.400 549.220 980.000 ;
      RECT 551.180 1.400 551.460 980.000 ;
      RECT 553.420 1.400 553.700 980.000 ;
      RECT 555.660 1.400 555.940 980.000 ;
      RECT 557.900 1.400 558.180 980.000 ;
      RECT 560.140 1.400 560.420 980.000 ;
      RECT 562.380 1.400 562.660 980.000 ;
      RECT 564.620 1.400 564.900 980.000 ;
      RECT 566.860 1.400 567.140 980.000 ;
      RECT 569.100 1.400 569.380 980.000 ;
      RECT 571.340 1.400 571.620 980.000 ;
      RECT 573.580 1.400 573.860 980.000 ;
      RECT 575.820 1.400 576.100 980.000 ;
      RECT 578.060 1.400 578.340 980.000 ;
      RECT 580.300 1.400 580.580 980.000 ;
      RECT 582.540 1.400 582.820 980.000 ;
      RECT 584.780 1.400 585.060 980.000 ;
      RECT 587.020 1.400 587.300 980.000 ;
      RECT 589.260 1.400 589.540 980.000 ;
      RECT 591.500 1.400 591.780 980.000 ;
      RECT 593.740 1.400 594.020 980.000 ;
      RECT 595.980 1.400 596.260 980.000 ;
      RECT 598.220 1.400 598.500 980.000 ;
      RECT 600.460 1.400 600.740 980.000 ;
      RECT 602.700 1.400 602.980 980.000 ;
      RECT 604.940 1.400 605.220 980.000 ;
      RECT 607.180 1.400 607.460 980.000 ;
      RECT 609.420 1.400 609.700 980.000 ;
      RECT 611.660 1.400 611.940 980.000 ;
      RECT 613.900 1.400 614.180 980.000 ;
      RECT 616.140 1.400 616.420 980.000 ;
      RECT 618.380 1.400 618.660 980.000 ;
      RECT 620.620 1.400 620.900 980.000 ;
      RECT 622.860 1.400 623.140 980.000 ;
      RECT 625.100 1.400 625.380 980.000 ;
      RECT 627.340 1.400 627.620 980.000 ;
      RECT 629.580 1.400 629.860 980.000 ;
      RECT 631.820 1.400 632.100 980.000 ;
      RECT 634.060 1.400 634.340 980.000 ;
      RECT 636.300 1.400 636.580 980.000 ;
      RECT 638.540 1.400 638.820 980.000 ;
      RECT 640.780 1.400 641.060 980.000 ;
      RECT 643.020 1.400 643.300 980.000 ;
      RECT 645.260 1.400 645.540 980.000 ;
      RECT 647.500 1.400 647.780 980.000 ;
      RECT 649.740 1.400 650.020 980.000 ;
      RECT 651.980 1.400 652.260 980.000 ;
      RECT 654.220 1.400 654.500 980.000 ;
      RECT 656.460 1.400 656.740 980.000 ;
      RECT 658.700 1.400 658.980 980.000 ;
      RECT 660.940 1.400 661.220 980.000 ;
      RECT 663.180 1.400 663.460 980.000 ;
      RECT 665.420 1.400 665.700 980.000 ;
      RECT 667.660 1.400 667.940 980.000 ;
      RECT 669.900 1.400 670.180 980.000 ;
      RECT 672.140 1.400 672.420 980.000 ;
      RECT 674.380 1.400 674.660 980.000 ;
      RECT 676.620 1.400 676.900 980.000 ;
      RECT 678.860 1.400 679.140 980.000 ;
      RECT 681.100 1.400 681.380 980.000 ;
      RECT 683.340 1.400 683.620 980.000 ;
      RECT 685.580 1.400 685.860 980.000 ;
      RECT 687.820 1.400 688.100 980.000 ;
      RECT 690.060 1.400 690.340 980.000 ;
      RECT 692.300 1.400 692.580 980.000 ;
      RECT 694.540 1.400 694.820 980.000 ;
      RECT 696.780 1.400 697.060 980.000 ;
      RECT 699.020 1.400 699.300 980.000 ;
      RECT 701.260 1.400 701.540 980.000 ;
      RECT 703.500 1.400 703.780 980.000 ;
      RECT 705.740 1.400 706.020 980.000 ;
      RECT 707.980 1.400 708.260 980.000 ;
      RECT 710.220 1.400 710.500 980.000 ;
      RECT 712.460 1.400 712.740 980.000 ;
      RECT 714.700 1.400 714.980 980.000 ;
      RECT 716.940 1.400 717.220 980.000 ;
      RECT 719.180 1.400 719.460 980.000 ;
      RECT 721.420 1.400 721.700 980.000 ;
      RECT 723.660 1.400 723.940 980.000 ;
      RECT 725.900 1.400 726.180 980.000 ;
      RECT 728.140 1.400 728.420 980.000 ;
      RECT 730.380 1.400 730.660 980.000 ;
      RECT 732.620 1.400 732.900 980.000 ;
      RECT 734.860 1.400 735.140 980.000 ;
      RECT 737.100 1.400 737.380 980.000 ;
      RECT 739.340 1.400 739.620 980.000 ;
      RECT 741.580 1.400 741.860 980.000 ;
      RECT 743.820 1.400 744.100 980.000 ;
      RECT 746.060 1.400 746.340 980.000 ;
      RECT 748.300 1.400 748.580 980.000 ;
      RECT 750.540 1.400 750.820 980.000 ;
      RECT 752.780 1.400 753.060 980.000 ;
      RECT 755.020 1.400 755.300 980.000 ;
      RECT 757.260 1.400 757.540 980.000 ;
      RECT 759.500 1.400 759.780 980.000 ;
      RECT 761.740 1.400 762.020 980.000 ;
      RECT 763.980 1.400 764.260 980.000 ;
      RECT 766.220 1.400 766.500 980.000 ;
      RECT 768.460 1.400 768.740 980.000 ;
      RECT 770.700 1.400 770.980 980.000 ;
      RECT 772.940 1.400 773.220 980.000 ;
      RECT 775.180 1.400 775.460 980.000 ;
      RECT 777.420 1.400 777.700 980.000 ;
      RECT 779.660 1.400 779.940 980.000 ;
      RECT 781.900 1.400 782.180 980.000 ;
      RECT 784.140 1.400 784.420 980.000 ;
      RECT 786.380 1.400 786.660 980.000 ;
      RECT 788.620 1.400 788.900 980.000 ;
      RECT 790.860 1.400 791.140 980.000 ;
      RECT 793.100 1.400 793.380 980.000 ;
      RECT 795.340 1.400 795.620 980.000 ;
      RECT 797.580 1.400 797.860 980.000 ;
      RECT 799.820 1.400 800.100 980.000 ;
      RECT 802.060 1.400 802.340 980.000 ;
      RECT 804.300 1.400 804.580 980.000 ;
      RECT 806.540 1.400 806.820 980.000 ;
      RECT 808.780 1.400 809.060 980.000 ;
      RECT 811.020 1.400 811.300 980.000 ;
      RECT 813.260 1.400 813.540 980.000 ;
      RECT 815.500 1.400 815.780 980.000 ;
      RECT 817.740 1.400 818.020 980.000 ;
      RECT 819.980 1.400 820.260 980.000 ;
      RECT 822.220 1.400 822.500 980.000 ;
      RECT 824.460 1.400 824.740 980.000 ;
      RECT 826.700 1.400 826.980 980.000 ;
      RECT 828.940 1.400 829.220 980.000 ;
      RECT 831.180 1.400 831.460 980.000 ;
      RECT 833.420 1.400 833.700 980.000 ;
      RECT 835.660 1.400 835.940 980.000 ;
      RECT 837.900 1.400 838.180 980.000 ;
      RECT 840.140 1.400 840.420 980.000 ;
      RECT 842.380 1.400 842.660 980.000 ;
      RECT 844.620 1.400 844.900 980.000 ;
      RECT 846.860 1.400 847.140 980.000 ;
      RECT 849.100 1.400 849.380 980.000 ;
      RECT 851.340 1.400 851.620 980.000 ;
      RECT 853.580 1.400 853.860 980.000 ;
      RECT 855.820 1.400 856.100 980.000 ;
      RECT 858.060 1.400 858.340 980.000 ;
      RECT 860.300 1.400 860.580 980.000 ;
      RECT 862.540 1.400 862.820 980.000 ;
      RECT 864.780 1.400 865.060 980.000 ;
      RECT 867.020 1.400 867.300 980.000 ;
      RECT 869.260 1.400 869.540 980.000 ;
      RECT 871.500 1.400 871.780 980.000 ;
      RECT 873.740 1.400 874.020 980.000 ;
      RECT 875.980 1.400 876.260 980.000 ;
      RECT 878.220 1.400 878.500 980.000 ;
      RECT 880.460 1.400 880.740 980.000 ;
      RECT 882.700 1.400 882.980 980.000 ;
      RECT 884.940 1.400 885.220 980.000 ;
      RECT 887.180 1.400 887.460 980.000 ;
      RECT 889.420 1.400 889.700 980.000 ;
      RECT 891.660 1.400 891.940 980.000 ;
      RECT 893.900 1.400 894.180 980.000 ;
      RECT 896.140 1.400 896.420 980.000 ;
      RECT 898.380 1.400 898.660 980.000 ;
      RECT 900.620 1.400 900.900 980.000 ;
      RECT 902.860 1.400 903.140 980.000 ;
      RECT 905.100 1.400 905.380 980.000 ;
      RECT 907.340 1.400 907.620 980.000 ;
      RECT 909.580 1.400 909.860 980.000 ;
      RECT 911.820 1.400 912.100 980.000 ;
      RECT 914.060 1.400 914.340 980.000 ;
      RECT 916.300 1.400 916.580 980.000 ;
      RECT 918.540 1.400 918.820 980.000 ;
      RECT 920.780 1.400 921.060 980.000 ;
      RECT 923.020 1.400 923.300 980.000 ;
      RECT 925.260 1.400 925.540 980.000 ;
      RECT 927.500 1.400 927.780 980.000 ;
      RECT 929.740 1.400 930.020 980.000 ;
      RECT 931.980 1.400 932.260 980.000 ;
      RECT 934.220 1.400 934.500 980.000 ;
      RECT 936.460 1.400 936.740 980.000 ;
      RECT 938.700 1.400 938.980 980.000 ;
      RECT 940.940 1.400 941.220 980.000 ;
      RECT 943.180 1.400 943.460 980.000 ;
      RECT 945.420 1.400 945.700 980.000 ;
      RECT 947.660 1.400 947.940 980.000 ;
      RECT 949.900 1.400 950.180 980.000 ;
      RECT 952.140 1.400 952.420 980.000 ;
      RECT 954.380 1.400 954.660 980.000 ;
      RECT 956.620 1.400 956.900 980.000 ;
      RECT 958.860 1.400 959.140 980.000 ;
      RECT 961.100 1.400 961.380 980.000 ;
      RECT 963.340 1.400 963.620 980.000 ;
      RECT 965.580 1.400 965.860 980.000 ;
      RECT 967.820 1.400 968.100 980.000 ;
      RECT 970.060 1.400 970.340 980.000 ;
      RECT 972.300 1.400 972.580 980.000 ;
      RECT 974.540 1.400 974.820 980.000 ;
      RECT 976.780 1.400 977.060 980.000 ;
      RECT 979.020 1.400 979.300 980.000 ;
      RECT 981.260 1.400 981.540 980.000 ;
      RECT 983.500 1.400 983.780 980.000 ;
      RECT 985.740 1.400 986.020 980.000 ;
      RECT 987.980 1.400 988.260 980.000 ;
      RECT 990.220 1.400 990.500 980.000 ;
      RECT 992.460 1.400 992.740 980.000 ;
      RECT 994.700 1.400 994.980 980.000 ;
      RECT 996.940 1.400 997.220 980.000 ;
      RECT 999.180 1.400 999.460 980.000 ;
      RECT 1001.420 1.400 1001.700 980.000 ;
      RECT 1003.660 1.400 1003.940 980.000 ;
      RECT 1005.900 1.400 1006.180 980.000 ;
      RECT 1008.140 1.400 1008.420 980.000 ;
      RECT 1010.380 1.400 1010.660 980.000 ;
      RECT 1012.620 1.400 1012.900 980.000 ;
      RECT 1014.860 1.400 1015.140 980.000 ;
      RECT 1017.100 1.400 1017.380 980.000 ;
      RECT 1019.340 1.400 1019.620 980.000 ;
      RECT 1021.580 1.400 1021.860 980.000 ;
      RECT 1023.820 1.400 1024.100 980.000 ;
      RECT 1026.060 1.400 1026.340 980.000 ;
      RECT 1028.300 1.400 1028.580 980.000 ;
      RECT 1030.540 1.400 1030.820 980.000 ;
      RECT 1032.780 1.400 1033.060 980.000 ;
      RECT 1035.020 1.400 1035.300 980.000 ;
      RECT 1037.260 1.400 1037.540 980.000 ;
      RECT 1039.500 1.400 1039.780 980.000 ;
      RECT 1041.740 1.400 1042.020 980.000 ;
      RECT 1043.980 1.400 1044.260 980.000 ;
      RECT 1046.220 1.400 1046.500 980.000 ;
      RECT 1048.460 1.400 1048.740 980.000 ;
      RECT 1050.700 1.400 1050.980 980.000 ;
      RECT 1052.940 1.400 1053.220 980.000 ;
      RECT 1055.180 1.400 1055.460 980.000 ;
      RECT 1057.420 1.400 1057.700 980.000 ;
      RECT 1059.660 1.400 1059.940 980.000 ;
      RECT 1061.900 1.400 1062.180 980.000 ;
      RECT 1064.140 1.400 1064.420 980.000 ;
      RECT 1066.380 1.400 1066.660 980.000 ;
      RECT 1068.620 1.400 1068.900 980.000 ;
      RECT 1070.860 1.400 1071.140 980.000 ;
      RECT 1073.100 1.400 1073.380 980.000 ;
      RECT 1075.340 1.400 1075.620 980.000 ;
      RECT 1077.580 1.400 1077.860 980.000 ;
      RECT 1079.820 1.400 1080.100 980.000 ;
      RECT 1082.060 1.400 1082.340 980.000 ;
      RECT 1084.300 1.400 1084.580 980.000 ;
      RECT 1086.540 1.400 1086.820 980.000 ;
      RECT 1088.780 1.400 1089.060 980.000 ;
      RECT 1091.020 1.400 1091.300 980.000 ;
      RECT 1093.260 1.400 1093.540 980.000 ;
      RECT 1095.500 1.400 1095.780 980.000 ;
      RECT 1097.740 1.400 1098.020 980.000 ;
      RECT 1099.980 1.400 1100.260 980.000 ;
      RECT 1102.220 1.400 1102.500 980.000 ;
      RECT 1104.460 1.400 1104.740 980.000 ;
      RECT 1106.700 1.400 1106.980 980.000 ;
      RECT 1108.940 1.400 1109.220 980.000 ;
      RECT 1111.180 1.400 1111.460 980.000 ;
      RECT 1113.420 1.400 1113.700 980.000 ;
      RECT 1115.660 1.400 1115.940 980.000 ;
      RECT 1117.900 1.400 1118.180 980.000 ;
      RECT 1120.140 1.400 1120.420 980.000 ;
      RECT 1122.380 1.400 1122.660 980.000 ;
      RECT 1124.620 1.400 1124.900 980.000 ;
      RECT 1126.860 1.400 1127.140 980.000 ;
      RECT 1129.100 1.400 1129.380 980.000 ;
      RECT 1131.340 1.400 1131.620 980.000 ;
      RECT 1133.580 1.400 1133.860 980.000 ;
      RECT 1135.820 1.400 1136.100 980.000 ;
      RECT 1138.060 1.400 1138.340 980.000 ;
      RECT 1140.300 1.400 1140.580 980.000 ;
      RECT 1142.540 1.400 1142.820 980.000 ;
      RECT 1144.780 1.400 1145.060 980.000 ;
      RECT 1147.020 1.400 1147.300 980.000 ;
      RECT 1149.260 1.400 1149.540 980.000 ;
      RECT 1151.500 1.400 1151.780 980.000 ;
      RECT 1153.740 1.400 1154.020 980.000 ;
      RECT 1155.980 1.400 1156.260 980.000 ;
      RECT 1158.220 1.400 1158.500 980.000 ;
      RECT 1160.460 1.400 1160.740 980.000 ;
      RECT 1162.700 1.400 1162.980 980.000 ;
      RECT 1164.940 1.400 1165.220 980.000 ;
      RECT 1167.180 1.400 1167.460 980.000 ;
      RECT 1169.420 1.400 1169.700 980.000 ;
      RECT 1171.660 1.400 1171.940 980.000 ;
      RECT 1173.900 1.400 1174.180 980.000 ;
      RECT 1176.140 1.400 1176.420 980.000 ;
      RECT 1178.380 1.400 1178.660 980.000 ;
      RECT 1180.620 1.400 1180.900 980.000 ;
      RECT 1182.860 1.400 1183.140 980.000 ;
      RECT 1185.100 1.400 1185.380 980.000 ;
      RECT 1187.340 1.400 1187.620 980.000 ;
      RECT 1189.580 1.400 1189.860 980.000 ;
      RECT 1191.820 1.400 1192.100 980.000 ;
      RECT 1194.060 1.400 1194.340 980.000 ;
      RECT 1196.300 1.400 1196.580 980.000 ;
      RECT 1198.540 1.400 1198.820 980.000 ;
      RECT 1200.780 1.400 1201.060 980.000 ;
      RECT 1203.020 1.400 1203.300 980.000 ;
      RECT 1205.260 1.400 1205.540 980.000 ;
      RECT 1207.500 1.400 1207.780 980.000 ;
      RECT 1209.740 1.400 1210.020 980.000 ;
      RECT 1211.980 1.400 1212.260 980.000 ;
      RECT 1214.220 1.400 1214.500 980.000 ;
      RECT 1216.460 1.400 1216.740 980.000 ;
      RECT 1218.700 1.400 1218.980 980.000 ;
      RECT 1220.940 1.400 1221.220 980.000 ;
      RECT 1223.180 1.400 1223.460 980.000 ;
      RECT 1225.420 1.400 1225.700 980.000 ;
      RECT 1227.660 1.400 1227.940 980.000 ;
      RECT 1229.900 1.400 1230.180 980.000 ;
      RECT 1232.140 1.400 1232.420 980.000 ;
      RECT 1234.380 1.400 1234.660 980.000 ;
      RECT 1236.620 1.400 1236.900 980.000 ;
      RECT 1238.860 1.400 1239.140 980.000 ;
      RECT 1241.100 1.400 1241.380 980.000 ;
      RECT 1243.340 1.400 1243.620 980.000 ;
      RECT 1245.580 1.400 1245.860 980.000 ;
      RECT 1247.820 1.400 1248.100 980.000 ;
      RECT 1250.060 1.400 1250.340 980.000 ;
      RECT 1252.300 1.400 1252.580 980.000 ;
      RECT 1254.540 1.400 1254.820 980.000 ;
      RECT 1256.780 1.400 1257.060 980.000 ;
      RECT 1259.020 1.400 1259.300 980.000 ;
      RECT 1261.260 1.400 1261.540 980.000 ;
      RECT 1263.500 1.400 1263.780 980.000 ;
      RECT 1265.740 1.400 1266.020 980.000 ;
      RECT 1267.980 1.400 1268.260 980.000 ;
      RECT 1270.220 1.400 1270.500 980.000 ;
      RECT 1272.460 1.400 1272.740 980.000 ;
      RECT 1274.700 1.400 1274.980 980.000 ;
      RECT 1276.940 1.400 1277.220 980.000 ;
      RECT 1279.180 1.400 1279.460 980.000 ;
      RECT 1281.420 1.400 1281.700 980.000 ;
      RECT 1283.660 1.400 1283.940 980.000 ;
      RECT 1285.900 1.400 1286.180 980.000 ;
      RECT 1288.140 1.400 1288.420 980.000 ;
      RECT 1290.380 1.400 1290.660 980.000 ;
      RECT 1292.620 1.400 1292.900 980.000 ;
      RECT 1294.860 1.400 1295.140 980.000 ;
      RECT 1297.100 1.400 1297.380 980.000 ;
      RECT 1299.340 1.400 1299.620 980.000 ;
      RECT 1301.580 1.400 1301.860 980.000 ;
      RECT 1303.820 1.400 1304.100 980.000 ;
      RECT 1306.060 1.400 1306.340 980.000 ;
      RECT 1308.300 1.400 1308.580 980.000 ;
      RECT 1310.540 1.400 1310.820 980.000 ;
      RECT 1312.780 1.400 1313.060 980.000 ;
      RECT 1315.020 1.400 1315.300 980.000 ;
      RECT 1317.260 1.400 1317.540 980.000 ;
      RECT 1319.500 1.400 1319.780 980.000 ;
      RECT 1321.740 1.400 1322.020 980.000 ;
      RECT 1323.980 1.400 1324.260 980.000 ;
      RECT 1326.220 1.400 1326.500 980.000 ;
      RECT 1328.460 1.400 1328.740 980.000 ;
      RECT 1330.700 1.400 1330.980 980.000 ;
      RECT 1332.940 1.400 1333.220 980.000 ;
      RECT 1335.180 1.400 1335.460 980.000 ;
      RECT 1337.420 1.400 1337.700 980.000 ;
      RECT 1339.660 1.400 1339.940 980.000 ;
      RECT 1341.900 1.400 1342.180 980.000 ;
      RECT 1344.140 1.400 1344.420 980.000 ;
      RECT 1346.380 1.400 1346.660 980.000 ;
      RECT 1348.620 1.400 1348.900 980.000 ;
      RECT 1350.860 1.400 1351.140 980.000 ;
      RECT 1353.100 1.400 1353.380 980.000 ;
      RECT 1355.340 1.400 1355.620 980.000 ;
      RECT 1357.580 1.400 1357.860 980.000 ;
      RECT 1359.820 1.400 1360.100 980.000 ;
      RECT 1362.060 1.400 1362.340 980.000 ;
      RECT 1364.300 1.400 1364.580 980.000 ;
      RECT 1366.540 1.400 1366.820 980.000 ;
      RECT 1368.780 1.400 1369.060 980.000 ;
      RECT 1371.020 1.400 1371.300 980.000 ;
      RECT 1373.260 1.400 1373.540 980.000 ;
      RECT 1375.500 1.400 1375.780 980.000 ;
      RECT 1377.740 1.400 1378.020 980.000 ;
      RECT 1379.980 1.400 1380.260 980.000 ;
      RECT 1382.220 1.400 1382.500 980.000 ;
      RECT 1384.460 1.400 1384.740 980.000 ;
      RECT 1386.700 1.400 1386.980 980.000 ;
      RECT 1388.940 1.400 1389.220 980.000 ;
      RECT 1391.180 1.400 1391.460 980.000 ;
      RECT 1393.420 1.400 1393.700 980.000 ;
      RECT 1395.660 1.400 1395.940 980.000 ;
      RECT 1397.900 1.400 1398.180 980.000 ;
      RECT 1400.140 1.400 1400.420 980.000 ;
      RECT 1402.380 1.400 1402.660 980.000 ;
      RECT 1404.620 1.400 1404.900 980.000 ;
      RECT 1406.860 1.400 1407.140 980.000 ;
      RECT 1409.100 1.400 1409.380 980.000 ;
      RECT 1411.340 1.400 1411.620 980.000 ;
      RECT 1413.580 1.400 1413.860 980.000 ;
      RECT 1415.820 1.400 1416.100 980.000 ;
      RECT 1418.060 1.400 1418.340 980.000 ;
      RECT 1420.300 1.400 1420.580 980.000 ;
      RECT 1422.540 1.400 1422.820 980.000 ;
      RECT 1424.780 1.400 1425.060 980.000 ;
      RECT 1427.020 1.400 1427.300 980.000 ;
      RECT 1429.260 1.400 1429.540 980.000 ;
      RECT 1431.500 1.400 1431.780 980.000 ;
      RECT 1433.740 1.400 1434.020 980.000 ;
      RECT 1435.980 1.400 1436.260 980.000 ;
      RECT 1438.220 1.400 1438.500 980.000 ;
      RECT 1440.460 1.400 1440.740 980.000 ;
      RECT 1442.700 1.400 1442.980 980.000 ;
      RECT 1444.940 1.400 1445.220 980.000 ;
      RECT 1447.180 1.400 1447.460 980.000 ;
      RECT 1449.420 1.400 1449.700 980.000 ;
      RECT 1451.660 1.400 1451.940 980.000 ;
      RECT 1453.900 1.400 1454.180 980.000 ;
      RECT 1456.140 1.400 1456.420 980.000 ;
      RECT 1458.380 1.400 1458.660 980.000 ;
      RECT 1460.620 1.400 1460.900 980.000 ;
      RECT 1462.860 1.400 1463.140 980.000 ;
      RECT 1465.100 1.400 1465.380 980.000 ;
      RECT 1467.340 1.400 1467.620 980.000 ;
      RECT 1469.580 1.400 1469.860 980.000 ;
      RECT 1471.820 1.400 1472.100 980.000 ;
      RECT 1474.060 1.400 1474.340 980.000 ;
      RECT 1476.300 1.400 1476.580 980.000 ;
      RECT 1478.540 1.400 1478.820 980.000 ;
      RECT 1480.780 1.400 1481.060 980.000 ;
      RECT 1483.020 1.400 1483.300 980.000 ;
      RECT 1485.260 1.400 1485.540 980.000 ;
      RECT 1487.500 1.400 1487.780 980.000 ;
      RECT 1489.740 1.400 1490.020 980.000 ;
      RECT 1491.980 1.400 1492.260 980.000 ;
      RECT 1494.220 1.400 1494.500 980.000 ;
      RECT 1496.460 1.400 1496.740 980.000 ;
      RECT 1498.700 1.400 1498.980 980.000 ;
      RECT 1500.940 1.400 1501.220 980.000 ;
      RECT 1503.180 1.400 1503.460 980.000 ;
      RECT 1505.420 1.400 1505.700 980.000 ;
      RECT 1507.660 1.400 1507.940 980.000 ;
      RECT 1509.900 1.400 1510.180 980.000 ;
      RECT 1512.140 1.400 1512.420 980.000 ;
      RECT 1514.380 1.400 1514.660 980.000 ;
      RECT 1516.620 1.400 1516.900 980.000 ;
      RECT 1518.860 1.400 1519.140 980.000 ;
      RECT 1521.100 1.400 1521.380 980.000 ;
      RECT 1523.340 1.400 1523.620 980.000 ;
      RECT 1525.580 1.400 1525.860 980.000 ;
      RECT 1527.820 1.400 1528.100 980.000 ;
      RECT 1530.060 1.400 1530.340 980.000 ;
      RECT 1532.300 1.400 1532.580 980.000 ;
      RECT 1534.540 1.400 1534.820 980.000 ;
      RECT 1536.780 1.400 1537.060 980.000 ;
      RECT 1539.020 1.400 1539.300 980.000 ;
      RECT 1541.260 1.400 1541.540 980.000 ;
      RECT 1543.500 1.400 1543.780 980.000 ;
      RECT 1545.740 1.400 1546.020 980.000 ;
      RECT 1547.980 1.400 1548.260 980.000 ;
      RECT 1550.220 1.400 1550.500 980.000 ;
      RECT 1552.460 1.400 1552.740 980.000 ;
      RECT 1554.700 1.400 1554.980 980.000 ;
      RECT 1556.940 1.400 1557.220 980.000 ;
      RECT 1559.180 1.400 1559.460 980.000 ;
      RECT 1561.420 1.400 1561.700 980.000 ;
      RECT 1563.660 1.400 1563.940 980.000 ;
      RECT 1565.900 1.400 1566.180 980.000 ;
      RECT 1568.140 1.400 1568.420 980.000 ;
      RECT 1570.380 1.400 1570.660 980.000 ;
      RECT 1572.620 1.400 1572.900 980.000 ;
      RECT 1574.860 1.400 1575.140 980.000 ;
      RECT 1577.100 1.400 1577.380 980.000 ;
      RECT 1579.340 1.400 1579.620 980.000 ;
      RECT 1581.580 1.400 1581.860 980.000 ;
      RECT 1583.820 1.400 1584.100 980.000 ;
      RECT 1586.060 1.400 1586.340 980.000 ;
      RECT 1588.300 1.400 1588.580 980.000 ;
      RECT 1590.540 1.400 1590.820 980.000 ;
      RECT 1592.780 1.400 1593.060 980.000 ;
      RECT 1595.020 1.400 1595.300 980.000 ;
      RECT 1597.260 1.400 1597.540 980.000 ;
      RECT 1599.500 1.400 1599.780 980.000 ;
      RECT 1601.740 1.400 1602.020 980.000 ;
      RECT 1603.980 1.400 1604.260 980.000 ;
      RECT 1606.220 1.400 1606.500 980.000 ;
      RECT 1608.460 1.400 1608.740 980.000 ;
      RECT 1610.700 1.400 1610.980 980.000 ;
      RECT 1612.940 1.400 1613.220 980.000 ;
      RECT 1615.180 1.400 1615.460 980.000 ;
      RECT 1617.420 1.400 1617.700 980.000 ;
      RECT 1619.660 1.400 1619.940 980.000 ;
      RECT 1621.900 1.400 1622.180 980.000 ;
      RECT 1624.140 1.400 1624.420 980.000 ;
      RECT 1626.380 1.400 1626.660 980.000 ;
      RECT 1628.620 1.400 1628.900 980.000 ;
      RECT 1630.860 1.400 1631.140 980.000 ;
      RECT 1633.100 1.400 1633.380 980.000 ;
      RECT 1635.340 1.400 1635.620 980.000 ;
      RECT 1637.580 1.400 1637.860 980.000 ;
      RECT 1639.820 1.400 1640.100 980.000 ;
      RECT 1642.060 1.400 1642.340 980.000 ;
      RECT 1644.300 1.400 1644.580 980.000 ;
      RECT 1646.540 1.400 1646.820 980.000 ;
      RECT 1648.780 1.400 1649.060 980.000 ;
      RECT 1651.020 1.400 1651.300 980.000 ;
      RECT 1653.260 1.400 1653.540 980.000 ;
      RECT 1655.500 1.400 1655.780 980.000 ;
      RECT 1657.740 1.400 1658.020 980.000 ;
      RECT 1659.980 1.400 1660.260 980.000 ;
      RECT 1662.220 1.400 1662.500 980.000 ;
      RECT 1664.460 1.400 1664.740 980.000 ;
      RECT 1666.700 1.400 1666.980 980.000 ;
      RECT 1668.940 1.400 1669.220 980.000 ;
      RECT 1671.180 1.400 1671.460 980.000 ;
      RECT 1673.420 1.400 1673.700 980.000 ;
      RECT 1675.660 1.400 1675.940 980.000 ;
      RECT 1677.900 1.400 1678.180 980.000 ;
      RECT 1680.140 1.400 1680.420 980.000 ;
      RECT 1682.380 1.400 1682.660 980.000 ;
      RECT 1684.620 1.400 1684.900 980.000 ;
      RECT 1686.860 1.400 1687.140 980.000 ;
      RECT 1689.100 1.400 1689.380 980.000 ;
      RECT 1691.340 1.400 1691.620 980.000 ;
      RECT 1693.580 1.400 1693.860 980.000 ;
      RECT 1695.820 1.400 1696.100 980.000 ;
      RECT 1698.060 1.400 1698.340 980.000 ;
      RECT 1700.300 1.400 1700.580 980.000 ;
      RECT 1702.540 1.400 1702.820 980.000 ;
      RECT 1704.780 1.400 1705.060 980.000 ;
      RECT 1707.020 1.400 1707.300 980.000 ;
      RECT 1709.260 1.400 1709.540 980.000 ;
      RECT 1711.500 1.400 1711.780 980.000 ;
      RECT 1713.740 1.400 1714.020 980.000 ;
      RECT 1715.980 1.400 1716.260 980.000 ;
      RECT 1718.220 1.400 1718.500 980.000 ;
      RECT 1720.460 1.400 1720.740 980.000 ;
      RECT 1722.700 1.400 1722.980 980.000 ;
      RECT 1724.940 1.400 1725.220 980.000 ;
      RECT 1727.180 1.400 1727.460 980.000 ;
      RECT 1729.420 1.400 1729.700 980.000 ;
      RECT 1731.660 1.400 1731.940 980.000 ;
      RECT 1733.900 1.400 1734.180 980.000 ;
      RECT 1736.140 1.400 1736.420 980.000 ;
      RECT 1738.380 1.400 1738.660 980.000 ;
      RECT 1740.620 1.400 1740.900 980.000 ;
      RECT 1742.860 1.400 1743.140 980.000 ;
      RECT 1745.100 1.400 1745.380 980.000 ;
      RECT 1747.340 1.400 1747.620 980.000 ;
      RECT 1749.580 1.400 1749.860 980.000 ;
      RECT 1751.820 1.400 1752.100 980.000 ;
      RECT 1754.060 1.400 1754.340 980.000 ;
      RECT 1756.300 1.400 1756.580 980.000 ;
      RECT 1758.540 1.400 1758.820 980.000 ;
      RECT 1760.780 1.400 1761.060 980.000 ;
      RECT 1763.020 1.400 1763.300 980.000 ;
      RECT 1765.260 1.400 1765.540 980.000 ;
      RECT 1767.500 1.400 1767.780 980.000 ;
      RECT 1769.740 1.400 1770.020 980.000 ;
      RECT 1771.980 1.400 1772.260 980.000 ;
      RECT 1774.220 1.400 1774.500 980.000 ;
      RECT 1776.460 1.400 1776.740 980.000 ;
      RECT 1778.700 1.400 1778.980 980.000 ;
      RECT 1780.940 1.400 1781.220 980.000 ;
      RECT 1783.180 1.400 1783.460 980.000 ;
      RECT 1785.420 1.400 1785.700 980.000 ;
      RECT 1787.660 1.400 1787.940 980.000 ;
      RECT 1789.900 1.400 1790.180 980.000 ;
      RECT 1792.140 1.400 1792.420 980.000 ;
      RECT 1794.380 1.400 1794.660 980.000 ;
      RECT 1796.620 1.400 1796.900 980.000 ;
      RECT 1798.860 1.400 1799.140 980.000 ;
      RECT 1801.100 1.400 1801.380 980.000 ;
      RECT 1803.340 1.400 1803.620 980.000 ;
      RECT 1805.580 1.400 1805.860 980.000 ;
      RECT 1807.820 1.400 1808.100 980.000 ;
      RECT 1810.060 1.400 1810.340 980.000 ;
      RECT 1812.300 1.400 1812.580 980.000 ;
      RECT 1814.540 1.400 1814.820 980.000 ;
      RECT 1816.780 1.400 1817.060 980.000 ;
      RECT 1819.020 1.400 1819.300 980.000 ;
      RECT 1821.260 1.400 1821.540 980.000 ;
      RECT 1823.500 1.400 1823.780 980.000 ;
      RECT 1825.740 1.400 1826.020 980.000 ;
      RECT 1827.980 1.400 1828.260 980.000 ;
      RECT 1830.220 1.400 1830.500 980.000 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 1832.740 981.400 ;
    LAYER metal2 ;
    RECT 0 0 1832.740 981.400 ;
    LAYER metal3 ;
    RECT 0.070 0 1832.740 981.400 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.925 ;
    RECT 0 1.995 0.070 2.485 ;
    RECT 0 2.555 0.070 3.045 ;
    RECT 0 3.115 0.070 3.605 ;
    RECT 0 3.675 0.070 4.165 ;
    RECT 0 4.235 0.070 4.725 ;
    RECT 0 4.795 0.070 5.285 ;
    RECT 0 5.355 0.070 5.845 ;
    RECT 0 5.915 0.070 6.405 ;
    RECT 0 6.475 0.070 6.965 ;
    RECT 0 7.035 0.070 7.525 ;
    RECT 0 7.595 0.070 8.085 ;
    RECT 0 8.155 0.070 8.645 ;
    RECT 0 8.715 0.070 9.205 ;
    RECT 0 9.275 0.070 9.765 ;
    RECT 0 9.835 0.070 10.325 ;
    RECT 0 10.395 0.070 10.885 ;
    RECT 0 10.955 0.070 11.445 ;
    RECT 0 11.515 0.070 12.005 ;
    RECT 0 12.075 0.070 12.565 ;
    RECT 0 12.635 0.070 13.125 ;
    RECT 0 13.195 0.070 13.685 ;
    RECT 0 13.755 0.070 14.245 ;
    RECT 0 14.315 0.070 14.805 ;
    RECT 0 14.875 0.070 15.365 ;
    RECT 0 15.435 0.070 15.925 ;
    RECT 0 15.995 0.070 16.485 ;
    RECT 0 16.555 0.070 17.045 ;
    RECT 0 17.115 0.070 17.605 ;
    RECT 0 17.675 0.070 18.165 ;
    RECT 0 18.235 0.070 18.725 ;
    RECT 0 18.795 0.070 19.285 ;
    RECT 0 19.355 0.070 19.845 ;
    RECT 0 19.915 0.070 20.405 ;
    RECT 0 20.475 0.070 20.965 ;
    RECT 0 21.035 0.070 21.525 ;
    RECT 0 21.595 0.070 22.085 ;
    RECT 0 22.155 0.070 22.645 ;
    RECT 0 22.715 0.070 23.205 ;
    RECT 0 23.275 0.070 23.765 ;
    RECT 0 23.835 0.070 24.325 ;
    RECT 0 24.395 0.070 24.885 ;
    RECT 0 24.955 0.070 25.445 ;
    RECT 0 25.515 0.070 26.005 ;
    RECT 0 26.075 0.070 26.565 ;
    RECT 0 26.635 0.070 27.125 ;
    RECT 0 27.195 0.070 27.685 ;
    RECT 0 27.755 0.070 28.245 ;
    RECT 0 28.315 0.070 28.805 ;
    RECT 0 28.875 0.070 29.365 ;
    RECT 0 29.435 0.070 29.925 ;
    RECT 0 29.995 0.070 30.485 ;
    RECT 0 30.555 0.070 31.045 ;
    RECT 0 31.115 0.070 31.605 ;
    RECT 0 31.675 0.070 32.165 ;
    RECT 0 32.235 0.070 32.725 ;
    RECT 0 32.795 0.070 33.285 ;
    RECT 0 33.355 0.070 33.845 ;
    RECT 0 33.915 0.070 34.405 ;
    RECT 0 34.475 0.070 34.965 ;
    RECT 0 35.035 0.070 35.525 ;
    RECT 0 35.595 0.070 36.085 ;
    RECT 0 36.155 0.070 36.645 ;
    RECT 0 36.715 0.070 37.205 ;
    RECT 0 37.275 0.070 37.765 ;
    RECT 0 37.835 0.070 38.325 ;
    RECT 0 38.395 0.070 38.885 ;
    RECT 0 38.955 0.070 39.445 ;
    RECT 0 39.515 0.070 40.005 ;
    RECT 0 40.075 0.070 40.565 ;
    RECT 0 40.635 0.070 41.125 ;
    RECT 0 41.195 0.070 41.685 ;
    RECT 0 41.755 0.070 42.245 ;
    RECT 0 42.315 0.070 42.805 ;
    RECT 0 42.875 0.070 43.365 ;
    RECT 0 43.435 0.070 43.925 ;
    RECT 0 43.995 0.070 44.485 ;
    RECT 0 44.555 0.070 45.045 ;
    RECT 0 45.115 0.070 45.605 ;
    RECT 0 45.675 0.070 46.165 ;
    RECT 0 46.235 0.070 46.725 ;
    RECT 0 46.795 0.070 47.285 ;
    RECT 0 47.355 0.070 47.845 ;
    RECT 0 47.915 0.070 48.405 ;
    RECT 0 48.475 0.070 48.965 ;
    RECT 0 49.035 0.070 49.525 ;
    RECT 0 49.595 0.070 50.085 ;
    RECT 0 50.155 0.070 50.645 ;
    RECT 0 50.715 0.070 51.205 ;
    RECT 0 51.275 0.070 51.765 ;
    RECT 0 51.835 0.070 52.325 ;
    RECT 0 52.395 0.070 52.885 ;
    RECT 0 52.955 0.070 53.445 ;
    RECT 0 53.515 0.070 54.005 ;
    RECT 0 54.075 0.070 54.565 ;
    RECT 0 54.635 0.070 55.125 ;
    RECT 0 55.195 0.070 55.685 ;
    RECT 0 55.755 0.070 56.245 ;
    RECT 0 56.315 0.070 56.805 ;
    RECT 0 56.875 0.070 57.365 ;
    RECT 0 57.435 0.070 57.925 ;
    RECT 0 57.995 0.070 58.485 ;
    RECT 0 58.555 0.070 59.045 ;
    RECT 0 59.115 0.070 59.605 ;
    RECT 0 59.675 0.070 60.165 ;
    RECT 0 60.235 0.070 60.725 ;
    RECT 0 60.795 0.070 61.285 ;
    RECT 0 61.355 0.070 61.845 ;
    RECT 0 61.915 0.070 62.405 ;
    RECT 0 62.475 0.070 62.965 ;
    RECT 0 63.035 0.070 63.525 ;
    RECT 0 63.595 0.070 64.085 ;
    RECT 0 64.155 0.070 64.645 ;
    RECT 0 64.715 0.070 65.205 ;
    RECT 0 65.275 0.070 65.765 ;
    RECT 0 65.835 0.070 66.325 ;
    RECT 0 66.395 0.070 66.885 ;
    RECT 0 66.955 0.070 67.445 ;
    RECT 0 67.515 0.070 68.005 ;
    RECT 0 68.075 0.070 68.565 ;
    RECT 0 68.635 0.070 69.125 ;
    RECT 0 69.195 0.070 69.685 ;
    RECT 0 69.755 0.070 70.245 ;
    RECT 0 70.315 0.070 70.805 ;
    RECT 0 70.875 0.070 71.365 ;
    RECT 0 71.435 0.070 71.925 ;
    RECT 0 71.995 0.070 72.485 ;
    RECT 0 72.555 0.070 73.045 ;
    RECT 0 73.115 0.070 73.605 ;
    RECT 0 73.675 0.070 74.165 ;
    RECT 0 74.235 0.070 74.725 ;
    RECT 0 74.795 0.070 75.285 ;
    RECT 0 75.355 0.070 75.845 ;
    RECT 0 75.915 0.070 76.405 ;
    RECT 0 76.475 0.070 76.965 ;
    RECT 0 77.035 0.070 77.525 ;
    RECT 0 77.595 0.070 78.085 ;
    RECT 0 78.155 0.070 78.645 ;
    RECT 0 78.715 0.070 79.205 ;
    RECT 0 79.275 0.070 79.765 ;
    RECT 0 79.835 0.070 80.325 ;
    RECT 0 80.395 0.070 80.885 ;
    RECT 0 80.955 0.070 81.445 ;
    RECT 0 81.515 0.070 82.005 ;
    RECT 0 82.075 0.070 82.565 ;
    RECT 0 82.635 0.070 83.125 ;
    RECT 0 83.195 0.070 83.685 ;
    RECT 0 83.755 0.070 84.245 ;
    RECT 0 84.315 0.070 84.805 ;
    RECT 0 84.875 0.070 85.365 ;
    RECT 0 85.435 0.070 85.925 ;
    RECT 0 85.995 0.070 86.485 ;
    RECT 0 86.555 0.070 87.045 ;
    RECT 0 87.115 0.070 87.605 ;
    RECT 0 87.675 0.070 88.165 ;
    RECT 0 88.235 0.070 88.725 ;
    RECT 0 88.795 0.070 89.285 ;
    RECT 0 89.355 0.070 89.845 ;
    RECT 0 89.915 0.070 90.405 ;
    RECT 0 90.475 0.070 90.965 ;
    RECT 0 91.035 0.070 91.525 ;
    RECT 0 91.595 0.070 92.085 ;
    RECT 0 92.155 0.070 92.645 ;
    RECT 0 92.715 0.070 93.205 ;
    RECT 0 93.275 0.070 93.765 ;
    RECT 0 93.835 0.070 94.325 ;
    RECT 0 94.395 0.070 94.885 ;
    RECT 0 94.955 0.070 95.445 ;
    RECT 0 95.515 0.070 96.005 ;
    RECT 0 96.075 0.070 96.565 ;
    RECT 0 96.635 0.070 97.125 ;
    RECT 0 97.195 0.070 97.685 ;
    RECT 0 97.755 0.070 98.245 ;
    RECT 0 98.315 0.070 98.805 ;
    RECT 0 98.875 0.070 99.365 ;
    RECT 0 99.435 0.070 99.925 ;
    RECT 0 99.995 0.070 100.485 ;
    RECT 0 100.555 0.070 101.045 ;
    RECT 0 101.115 0.070 101.605 ;
    RECT 0 101.675 0.070 102.165 ;
    RECT 0 102.235 0.070 102.725 ;
    RECT 0 102.795 0.070 103.285 ;
    RECT 0 103.355 0.070 103.845 ;
    RECT 0 103.915 0.070 104.405 ;
    RECT 0 104.475 0.070 104.965 ;
    RECT 0 105.035 0.070 105.525 ;
    RECT 0 105.595 0.070 106.085 ;
    RECT 0 106.155 0.070 106.645 ;
    RECT 0 106.715 0.070 107.205 ;
    RECT 0 107.275 0.070 107.765 ;
    RECT 0 107.835 0.070 108.325 ;
    RECT 0 108.395 0.070 108.885 ;
    RECT 0 108.955 0.070 109.445 ;
    RECT 0 109.515 0.070 110.005 ;
    RECT 0 110.075 0.070 110.565 ;
    RECT 0 110.635 0.070 111.125 ;
    RECT 0 111.195 0.070 111.685 ;
    RECT 0 111.755 0.070 112.245 ;
    RECT 0 112.315 0.070 112.805 ;
    RECT 0 112.875 0.070 113.365 ;
    RECT 0 113.435 0.070 113.925 ;
    RECT 0 113.995 0.070 114.485 ;
    RECT 0 114.555 0.070 115.045 ;
    RECT 0 115.115 0.070 115.605 ;
    RECT 0 115.675 0.070 116.165 ;
    RECT 0 116.235 0.070 116.725 ;
    RECT 0 116.795 0.070 117.285 ;
    RECT 0 117.355 0.070 117.845 ;
    RECT 0 117.915 0.070 118.405 ;
    RECT 0 118.475 0.070 118.965 ;
    RECT 0 119.035 0.070 119.525 ;
    RECT 0 119.595 0.070 120.085 ;
    RECT 0 120.155 0.070 120.645 ;
    RECT 0 120.715 0.070 121.205 ;
    RECT 0 121.275 0.070 121.765 ;
    RECT 0 121.835 0.070 122.325 ;
    RECT 0 122.395 0.070 122.885 ;
    RECT 0 122.955 0.070 123.445 ;
    RECT 0 123.515 0.070 124.005 ;
    RECT 0 124.075 0.070 124.565 ;
    RECT 0 124.635 0.070 125.125 ;
    RECT 0 125.195 0.070 125.685 ;
    RECT 0 125.755 0.070 126.245 ;
    RECT 0 126.315 0.070 126.805 ;
    RECT 0 126.875 0.070 127.365 ;
    RECT 0 127.435 0.070 127.925 ;
    RECT 0 127.995 0.070 128.485 ;
    RECT 0 128.555 0.070 129.045 ;
    RECT 0 129.115 0.070 129.605 ;
    RECT 0 129.675 0.070 130.165 ;
    RECT 0 130.235 0.070 130.725 ;
    RECT 0 130.795 0.070 131.285 ;
    RECT 0 131.355 0.070 131.845 ;
    RECT 0 131.915 0.070 132.405 ;
    RECT 0 132.475 0.070 132.965 ;
    RECT 0 133.035 0.070 133.525 ;
    RECT 0 133.595 0.070 134.085 ;
    RECT 0 134.155 0.070 134.645 ;
    RECT 0 134.715 0.070 135.205 ;
    RECT 0 135.275 0.070 135.765 ;
    RECT 0 135.835 0.070 136.325 ;
    RECT 0 136.395 0.070 136.885 ;
    RECT 0 136.955 0.070 137.445 ;
    RECT 0 137.515 0.070 138.005 ;
    RECT 0 138.075 0.070 138.565 ;
    RECT 0 138.635 0.070 139.125 ;
    RECT 0 139.195 0.070 139.685 ;
    RECT 0 139.755 0.070 140.245 ;
    RECT 0 140.315 0.070 140.805 ;
    RECT 0 140.875 0.070 141.365 ;
    RECT 0 141.435 0.070 141.925 ;
    RECT 0 141.995 0.070 142.485 ;
    RECT 0 142.555 0.070 143.045 ;
    RECT 0 143.115 0.070 143.605 ;
    RECT 0 143.675 0.070 144.165 ;
    RECT 0 144.235 0.070 144.725 ;
    RECT 0 144.795 0.070 145.285 ;
    RECT 0 145.355 0.070 145.845 ;
    RECT 0 145.915 0.070 146.405 ;
    RECT 0 146.475 0.070 146.965 ;
    RECT 0 147.035 0.070 147.525 ;
    RECT 0 147.595 0.070 148.085 ;
    RECT 0 148.155 0.070 148.645 ;
    RECT 0 148.715 0.070 149.205 ;
    RECT 0 149.275 0.070 149.765 ;
    RECT 0 149.835 0.070 150.325 ;
    RECT 0 150.395 0.070 150.885 ;
    RECT 0 150.955 0.070 151.445 ;
    RECT 0 151.515 0.070 152.005 ;
    RECT 0 152.075 0.070 152.565 ;
    RECT 0 152.635 0.070 153.125 ;
    RECT 0 153.195 0.070 153.685 ;
    RECT 0 153.755 0.070 154.245 ;
    RECT 0 154.315 0.070 154.805 ;
    RECT 0 154.875 0.070 155.365 ;
    RECT 0 155.435 0.070 155.925 ;
    RECT 0 155.995 0.070 156.485 ;
    RECT 0 156.555 0.070 157.045 ;
    RECT 0 157.115 0.070 157.605 ;
    RECT 0 157.675 0.070 158.165 ;
    RECT 0 158.235 0.070 158.725 ;
    RECT 0 158.795 0.070 159.285 ;
    RECT 0 159.355 0.070 159.845 ;
    RECT 0 159.915 0.070 160.405 ;
    RECT 0 160.475 0.070 160.965 ;
    RECT 0 161.035 0.070 161.525 ;
    RECT 0 161.595 0.070 162.085 ;
    RECT 0 162.155 0.070 162.645 ;
    RECT 0 162.715 0.070 163.205 ;
    RECT 0 163.275 0.070 163.765 ;
    RECT 0 163.835 0.070 164.325 ;
    RECT 0 164.395 0.070 164.885 ;
    RECT 0 164.955 0.070 165.445 ;
    RECT 0 165.515 0.070 166.005 ;
    RECT 0 166.075 0.070 166.565 ;
    RECT 0 166.635 0.070 167.125 ;
    RECT 0 167.195 0.070 167.685 ;
    RECT 0 167.755 0.070 168.245 ;
    RECT 0 168.315 0.070 168.805 ;
    RECT 0 168.875 0.070 169.365 ;
    RECT 0 169.435 0.070 169.925 ;
    RECT 0 169.995 0.070 170.485 ;
    RECT 0 170.555 0.070 171.045 ;
    RECT 0 171.115 0.070 171.605 ;
    RECT 0 171.675 0.070 172.165 ;
    RECT 0 172.235 0.070 172.725 ;
    RECT 0 172.795 0.070 173.285 ;
    RECT 0 173.355 0.070 173.845 ;
    RECT 0 173.915 0.070 174.405 ;
    RECT 0 174.475 0.070 174.965 ;
    RECT 0 175.035 0.070 175.525 ;
    RECT 0 175.595 0.070 176.085 ;
    RECT 0 176.155 0.070 176.645 ;
    RECT 0 176.715 0.070 177.205 ;
    RECT 0 177.275 0.070 177.765 ;
    RECT 0 177.835 0.070 178.325 ;
    RECT 0 178.395 0.070 178.885 ;
    RECT 0 178.955 0.070 179.445 ;
    RECT 0 179.515 0.070 180.005 ;
    RECT 0 180.075 0.070 180.565 ;
    RECT 0 180.635 0.070 181.125 ;
    RECT 0 181.195 0.070 181.685 ;
    RECT 0 181.755 0.070 182.245 ;
    RECT 0 182.315 0.070 182.805 ;
    RECT 0 182.875 0.070 183.365 ;
    RECT 0 183.435 0.070 183.925 ;
    RECT 0 183.995 0.070 184.485 ;
    RECT 0 184.555 0.070 185.045 ;
    RECT 0 185.115 0.070 185.605 ;
    RECT 0 185.675 0.070 186.165 ;
    RECT 0 186.235 0.070 186.725 ;
    RECT 0 186.795 0.070 187.285 ;
    RECT 0 187.355 0.070 187.845 ;
    RECT 0 187.915 0.070 188.405 ;
    RECT 0 188.475 0.070 188.965 ;
    RECT 0 189.035 0.070 189.525 ;
    RECT 0 189.595 0.070 190.085 ;
    RECT 0 190.155 0.070 190.645 ;
    RECT 0 190.715 0.070 191.205 ;
    RECT 0 191.275 0.070 191.765 ;
    RECT 0 191.835 0.070 192.325 ;
    RECT 0 192.395 0.070 192.885 ;
    RECT 0 192.955 0.070 193.445 ;
    RECT 0 193.515 0.070 194.005 ;
    RECT 0 194.075 0.070 194.565 ;
    RECT 0 194.635 0.070 195.125 ;
    RECT 0 195.195 0.070 195.685 ;
    RECT 0 195.755 0.070 196.245 ;
    RECT 0 196.315 0.070 196.805 ;
    RECT 0 196.875 0.070 197.365 ;
    RECT 0 197.435 0.070 197.925 ;
    RECT 0 197.995 0.070 198.485 ;
    RECT 0 198.555 0.070 199.045 ;
    RECT 0 199.115 0.070 199.605 ;
    RECT 0 199.675 0.070 200.165 ;
    RECT 0 200.235 0.070 200.725 ;
    RECT 0 200.795 0.070 201.285 ;
    RECT 0 201.355 0.070 201.845 ;
    RECT 0 201.915 0.070 202.405 ;
    RECT 0 202.475 0.070 202.965 ;
    RECT 0 203.035 0.070 203.525 ;
    RECT 0 203.595 0.070 204.085 ;
    RECT 0 204.155 0.070 204.645 ;
    RECT 0 204.715 0.070 205.205 ;
    RECT 0 205.275 0.070 205.765 ;
    RECT 0 205.835 0.070 206.325 ;
    RECT 0 206.395 0.070 206.885 ;
    RECT 0 206.955 0.070 207.445 ;
    RECT 0 207.515 0.070 208.005 ;
    RECT 0 208.075 0.070 208.565 ;
    RECT 0 208.635 0.070 209.125 ;
    RECT 0 209.195 0.070 209.685 ;
    RECT 0 209.755 0.070 210.245 ;
    RECT 0 210.315 0.070 210.805 ;
    RECT 0 210.875 0.070 211.365 ;
    RECT 0 211.435 0.070 211.925 ;
    RECT 0 211.995 0.070 212.485 ;
    RECT 0 212.555 0.070 213.045 ;
    RECT 0 213.115 0.070 213.605 ;
    RECT 0 213.675 0.070 214.165 ;
    RECT 0 214.235 0.070 214.725 ;
    RECT 0 214.795 0.070 215.285 ;
    RECT 0 215.355 0.070 215.845 ;
    RECT 0 215.915 0.070 216.405 ;
    RECT 0 216.475 0.070 216.965 ;
    RECT 0 217.035 0.070 217.525 ;
    RECT 0 217.595 0.070 218.085 ;
    RECT 0 218.155 0.070 218.645 ;
    RECT 0 218.715 0.070 219.205 ;
    RECT 0 219.275 0.070 219.765 ;
    RECT 0 219.835 0.070 220.325 ;
    RECT 0 220.395 0.070 220.885 ;
    RECT 0 220.955 0.070 221.445 ;
    RECT 0 221.515 0.070 222.005 ;
    RECT 0 222.075 0.070 222.565 ;
    RECT 0 222.635 0.070 223.125 ;
    RECT 0 223.195 0.070 223.685 ;
    RECT 0 223.755 0.070 224.245 ;
    RECT 0 224.315 0.070 224.805 ;
    RECT 0 224.875 0.070 225.365 ;
    RECT 0 225.435 0.070 225.925 ;
    RECT 0 225.995 0.070 226.485 ;
    RECT 0 226.555 0.070 227.045 ;
    RECT 0 227.115 0.070 227.605 ;
    RECT 0 227.675 0.070 228.165 ;
    RECT 0 228.235 0.070 228.725 ;
    RECT 0 228.795 0.070 229.285 ;
    RECT 0 229.355 0.070 229.845 ;
    RECT 0 229.915 0.070 230.405 ;
    RECT 0 230.475 0.070 230.965 ;
    RECT 0 231.035 0.070 231.525 ;
    RECT 0 231.595 0.070 232.085 ;
    RECT 0 232.155 0.070 232.645 ;
    RECT 0 232.715 0.070 233.205 ;
    RECT 0 233.275 0.070 233.765 ;
    RECT 0 233.835 0.070 234.325 ;
    RECT 0 234.395 0.070 234.885 ;
    RECT 0 234.955 0.070 235.445 ;
    RECT 0 235.515 0.070 236.005 ;
    RECT 0 236.075 0.070 236.565 ;
    RECT 0 236.635 0.070 237.125 ;
    RECT 0 237.195 0.070 237.685 ;
    RECT 0 237.755 0.070 238.245 ;
    RECT 0 238.315 0.070 238.805 ;
    RECT 0 238.875 0.070 239.365 ;
    RECT 0 239.435 0.070 239.925 ;
    RECT 0 239.995 0.070 240.485 ;
    RECT 0 240.555 0.070 241.045 ;
    RECT 0 241.115 0.070 241.605 ;
    RECT 0 241.675 0.070 242.165 ;
    RECT 0 242.235 0.070 242.725 ;
    RECT 0 242.795 0.070 243.285 ;
    RECT 0 243.355 0.070 243.845 ;
    RECT 0 243.915 0.070 244.405 ;
    RECT 0 244.475 0.070 244.965 ;
    RECT 0 245.035 0.070 245.525 ;
    RECT 0 245.595 0.070 246.085 ;
    RECT 0 246.155 0.070 246.645 ;
    RECT 0 246.715 0.070 247.205 ;
    RECT 0 247.275 0.070 247.765 ;
    RECT 0 247.835 0.070 248.325 ;
    RECT 0 248.395 0.070 248.885 ;
    RECT 0 248.955 0.070 249.445 ;
    RECT 0 249.515 0.070 250.005 ;
    RECT 0 250.075 0.070 250.565 ;
    RECT 0 250.635 0.070 251.125 ;
    RECT 0 251.195 0.070 251.685 ;
    RECT 0 251.755 0.070 252.245 ;
    RECT 0 252.315 0.070 252.805 ;
    RECT 0 252.875 0.070 253.365 ;
    RECT 0 253.435 0.070 253.925 ;
    RECT 0 253.995 0.070 254.485 ;
    RECT 0 254.555 0.070 255.045 ;
    RECT 0 255.115 0.070 255.605 ;
    RECT 0 255.675 0.070 256.165 ;
    RECT 0 256.235 0.070 256.725 ;
    RECT 0 256.795 0.070 257.285 ;
    RECT 0 257.355 0.070 257.845 ;
    RECT 0 257.915 0.070 258.405 ;
    RECT 0 258.475 0.070 258.965 ;
    RECT 0 259.035 0.070 259.525 ;
    RECT 0 259.595 0.070 260.085 ;
    RECT 0 260.155 0.070 260.645 ;
    RECT 0 260.715 0.070 261.205 ;
    RECT 0 261.275 0.070 261.765 ;
    RECT 0 261.835 0.070 262.325 ;
    RECT 0 262.395 0.070 262.885 ;
    RECT 0 262.955 0.070 263.445 ;
    RECT 0 263.515 0.070 264.005 ;
    RECT 0 264.075 0.070 264.565 ;
    RECT 0 264.635 0.070 265.125 ;
    RECT 0 265.195 0.070 265.685 ;
    RECT 0 265.755 0.070 266.245 ;
    RECT 0 266.315 0.070 266.805 ;
    RECT 0 266.875 0.070 267.365 ;
    RECT 0 267.435 0.070 267.925 ;
    RECT 0 267.995 0.070 268.485 ;
    RECT 0 268.555 0.070 269.045 ;
    RECT 0 269.115 0.070 269.605 ;
    RECT 0 269.675 0.070 270.165 ;
    RECT 0 270.235 0.070 270.725 ;
    RECT 0 270.795 0.070 271.285 ;
    RECT 0 271.355 0.070 271.845 ;
    RECT 0 271.915 0.070 272.405 ;
    RECT 0 272.475 0.070 272.965 ;
    RECT 0 273.035 0.070 273.525 ;
    RECT 0 273.595 0.070 274.085 ;
    RECT 0 274.155 0.070 274.645 ;
    RECT 0 274.715 0.070 275.205 ;
    RECT 0 275.275 0.070 275.765 ;
    RECT 0 275.835 0.070 276.325 ;
    RECT 0 276.395 0.070 276.885 ;
    RECT 0 276.955 0.070 277.445 ;
    RECT 0 277.515 0.070 278.005 ;
    RECT 0 278.075 0.070 278.565 ;
    RECT 0 278.635 0.070 279.125 ;
    RECT 0 279.195 0.070 279.685 ;
    RECT 0 279.755 0.070 280.245 ;
    RECT 0 280.315 0.070 280.805 ;
    RECT 0 280.875 0.070 281.365 ;
    RECT 0 281.435 0.070 281.925 ;
    RECT 0 281.995 0.070 282.485 ;
    RECT 0 282.555 0.070 283.045 ;
    RECT 0 283.115 0.070 283.605 ;
    RECT 0 283.675 0.070 284.165 ;
    RECT 0 284.235 0.070 284.725 ;
    RECT 0 284.795 0.070 285.285 ;
    RECT 0 285.355 0.070 285.845 ;
    RECT 0 285.915 0.070 286.405 ;
    RECT 0 286.475 0.070 286.965 ;
    RECT 0 287.035 0.070 287.525 ;
    RECT 0 287.595 0.070 315.245 ;
    RECT 0 315.315 0.070 315.805 ;
    RECT 0 315.875 0.070 316.365 ;
    RECT 0 316.435 0.070 316.925 ;
    RECT 0 316.995 0.070 317.485 ;
    RECT 0 317.555 0.070 318.045 ;
    RECT 0 318.115 0.070 318.605 ;
    RECT 0 318.675 0.070 319.165 ;
    RECT 0 319.235 0.070 319.725 ;
    RECT 0 319.795 0.070 320.285 ;
    RECT 0 320.355 0.070 320.845 ;
    RECT 0 320.915 0.070 321.405 ;
    RECT 0 321.475 0.070 321.965 ;
    RECT 0 322.035 0.070 322.525 ;
    RECT 0 322.595 0.070 323.085 ;
    RECT 0 323.155 0.070 323.645 ;
    RECT 0 323.715 0.070 324.205 ;
    RECT 0 324.275 0.070 324.765 ;
    RECT 0 324.835 0.070 325.325 ;
    RECT 0 325.395 0.070 325.885 ;
    RECT 0 325.955 0.070 326.445 ;
    RECT 0 326.515 0.070 327.005 ;
    RECT 0 327.075 0.070 327.565 ;
    RECT 0 327.635 0.070 328.125 ;
    RECT 0 328.195 0.070 328.685 ;
    RECT 0 328.755 0.070 329.245 ;
    RECT 0 329.315 0.070 329.805 ;
    RECT 0 329.875 0.070 330.365 ;
    RECT 0 330.435 0.070 330.925 ;
    RECT 0 330.995 0.070 331.485 ;
    RECT 0 331.555 0.070 332.045 ;
    RECT 0 332.115 0.070 332.605 ;
    RECT 0 332.675 0.070 333.165 ;
    RECT 0 333.235 0.070 333.725 ;
    RECT 0 333.795 0.070 334.285 ;
    RECT 0 334.355 0.070 334.845 ;
    RECT 0 334.915 0.070 335.405 ;
    RECT 0 335.475 0.070 335.965 ;
    RECT 0 336.035 0.070 336.525 ;
    RECT 0 336.595 0.070 337.085 ;
    RECT 0 337.155 0.070 337.645 ;
    RECT 0 337.715 0.070 338.205 ;
    RECT 0 338.275 0.070 338.765 ;
    RECT 0 338.835 0.070 339.325 ;
    RECT 0 339.395 0.070 339.885 ;
    RECT 0 339.955 0.070 340.445 ;
    RECT 0 340.515 0.070 341.005 ;
    RECT 0 341.075 0.070 341.565 ;
    RECT 0 341.635 0.070 342.125 ;
    RECT 0 342.195 0.070 342.685 ;
    RECT 0 342.755 0.070 343.245 ;
    RECT 0 343.315 0.070 343.805 ;
    RECT 0 343.875 0.070 344.365 ;
    RECT 0 344.435 0.070 344.925 ;
    RECT 0 344.995 0.070 345.485 ;
    RECT 0 345.555 0.070 346.045 ;
    RECT 0 346.115 0.070 346.605 ;
    RECT 0 346.675 0.070 347.165 ;
    RECT 0 347.235 0.070 347.725 ;
    RECT 0 347.795 0.070 348.285 ;
    RECT 0 348.355 0.070 348.845 ;
    RECT 0 348.915 0.070 349.405 ;
    RECT 0 349.475 0.070 349.965 ;
    RECT 0 350.035 0.070 350.525 ;
    RECT 0 350.595 0.070 351.085 ;
    RECT 0 351.155 0.070 351.645 ;
    RECT 0 351.715 0.070 352.205 ;
    RECT 0 352.275 0.070 352.765 ;
    RECT 0 352.835 0.070 353.325 ;
    RECT 0 353.395 0.070 353.885 ;
    RECT 0 353.955 0.070 354.445 ;
    RECT 0 354.515 0.070 355.005 ;
    RECT 0 355.075 0.070 355.565 ;
    RECT 0 355.635 0.070 356.125 ;
    RECT 0 356.195 0.070 356.685 ;
    RECT 0 356.755 0.070 357.245 ;
    RECT 0 357.315 0.070 357.805 ;
    RECT 0 357.875 0.070 358.365 ;
    RECT 0 358.435 0.070 358.925 ;
    RECT 0 358.995 0.070 359.485 ;
    RECT 0 359.555 0.070 360.045 ;
    RECT 0 360.115 0.070 360.605 ;
    RECT 0 360.675 0.070 361.165 ;
    RECT 0 361.235 0.070 361.725 ;
    RECT 0 361.795 0.070 362.285 ;
    RECT 0 362.355 0.070 362.845 ;
    RECT 0 362.915 0.070 363.405 ;
    RECT 0 363.475 0.070 363.965 ;
    RECT 0 364.035 0.070 364.525 ;
    RECT 0 364.595 0.070 365.085 ;
    RECT 0 365.155 0.070 365.645 ;
    RECT 0 365.715 0.070 366.205 ;
    RECT 0 366.275 0.070 366.765 ;
    RECT 0 366.835 0.070 367.325 ;
    RECT 0 367.395 0.070 367.885 ;
    RECT 0 367.955 0.070 368.445 ;
    RECT 0 368.515 0.070 369.005 ;
    RECT 0 369.075 0.070 369.565 ;
    RECT 0 369.635 0.070 370.125 ;
    RECT 0 370.195 0.070 370.685 ;
    RECT 0 370.755 0.070 371.245 ;
    RECT 0 371.315 0.070 371.805 ;
    RECT 0 371.875 0.070 372.365 ;
    RECT 0 372.435 0.070 372.925 ;
    RECT 0 372.995 0.070 373.485 ;
    RECT 0 373.555 0.070 374.045 ;
    RECT 0 374.115 0.070 374.605 ;
    RECT 0 374.675 0.070 375.165 ;
    RECT 0 375.235 0.070 375.725 ;
    RECT 0 375.795 0.070 376.285 ;
    RECT 0 376.355 0.070 376.845 ;
    RECT 0 376.915 0.070 377.405 ;
    RECT 0 377.475 0.070 377.965 ;
    RECT 0 378.035 0.070 378.525 ;
    RECT 0 378.595 0.070 379.085 ;
    RECT 0 379.155 0.070 379.645 ;
    RECT 0 379.715 0.070 380.205 ;
    RECT 0 380.275 0.070 380.765 ;
    RECT 0 380.835 0.070 381.325 ;
    RECT 0 381.395 0.070 381.885 ;
    RECT 0 381.955 0.070 382.445 ;
    RECT 0 382.515 0.070 383.005 ;
    RECT 0 383.075 0.070 383.565 ;
    RECT 0 383.635 0.070 384.125 ;
    RECT 0 384.195 0.070 384.685 ;
    RECT 0 384.755 0.070 385.245 ;
    RECT 0 385.315 0.070 385.805 ;
    RECT 0 385.875 0.070 386.365 ;
    RECT 0 386.435 0.070 386.925 ;
    RECT 0 386.995 0.070 387.485 ;
    RECT 0 387.555 0.070 388.045 ;
    RECT 0 388.115 0.070 388.605 ;
    RECT 0 388.675 0.070 389.165 ;
    RECT 0 389.235 0.070 389.725 ;
    RECT 0 389.795 0.070 390.285 ;
    RECT 0 390.355 0.070 390.845 ;
    RECT 0 390.915 0.070 391.405 ;
    RECT 0 391.475 0.070 391.965 ;
    RECT 0 392.035 0.070 392.525 ;
    RECT 0 392.595 0.070 393.085 ;
    RECT 0 393.155 0.070 393.645 ;
    RECT 0 393.715 0.070 394.205 ;
    RECT 0 394.275 0.070 394.765 ;
    RECT 0 394.835 0.070 395.325 ;
    RECT 0 395.395 0.070 395.885 ;
    RECT 0 395.955 0.070 396.445 ;
    RECT 0 396.515 0.070 397.005 ;
    RECT 0 397.075 0.070 397.565 ;
    RECT 0 397.635 0.070 398.125 ;
    RECT 0 398.195 0.070 398.685 ;
    RECT 0 398.755 0.070 399.245 ;
    RECT 0 399.315 0.070 399.805 ;
    RECT 0 399.875 0.070 400.365 ;
    RECT 0 400.435 0.070 400.925 ;
    RECT 0 400.995 0.070 401.485 ;
    RECT 0 401.555 0.070 402.045 ;
    RECT 0 402.115 0.070 402.605 ;
    RECT 0 402.675 0.070 403.165 ;
    RECT 0 403.235 0.070 403.725 ;
    RECT 0 403.795 0.070 404.285 ;
    RECT 0 404.355 0.070 404.845 ;
    RECT 0 404.915 0.070 405.405 ;
    RECT 0 405.475 0.070 405.965 ;
    RECT 0 406.035 0.070 406.525 ;
    RECT 0 406.595 0.070 407.085 ;
    RECT 0 407.155 0.070 407.645 ;
    RECT 0 407.715 0.070 408.205 ;
    RECT 0 408.275 0.070 408.765 ;
    RECT 0 408.835 0.070 409.325 ;
    RECT 0 409.395 0.070 409.885 ;
    RECT 0 409.955 0.070 410.445 ;
    RECT 0 410.515 0.070 411.005 ;
    RECT 0 411.075 0.070 411.565 ;
    RECT 0 411.635 0.070 412.125 ;
    RECT 0 412.195 0.070 412.685 ;
    RECT 0 412.755 0.070 413.245 ;
    RECT 0 413.315 0.070 413.805 ;
    RECT 0 413.875 0.070 414.365 ;
    RECT 0 414.435 0.070 414.925 ;
    RECT 0 414.995 0.070 415.485 ;
    RECT 0 415.555 0.070 416.045 ;
    RECT 0 416.115 0.070 416.605 ;
    RECT 0 416.675 0.070 417.165 ;
    RECT 0 417.235 0.070 417.725 ;
    RECT 0 417.795 0.070 418.285 ;
    RECT 0 418.355 0.070 418.845 ;
    RECT 0 418.915 0.070 419.405 ;
    RECT 0 419.475 0.070 419.965 ;
    RECT 0 420.035 0.070 420.525 ;
    RECT 0 420.595 0.070 421.085 ;
    RECT 0 421.155 0.070 421.645 ;
    RECT 0 421.715 0.070 422.205 ;
    RECT 0 422.275 0.070 422.765 ;
    RECT 0 422.835 0.070 423.325 ;
    RECT 0 423.395 0.070 423.885 ;
    RECT 0 423.955 0.070 424.445 ;
    RECT 0 424.515 0.070 425.005 ;
    RECT 0 425.075 0.070 425.565 ;
    RECT 0 425.635 0.070 426.125 ;
    RECT 0 426.195 0.070 426.685 ;
    RECT 0 426.755 0.070 427.245 ;
    RECT 0 427.315 0.070 427.805 ;
    RECT 0 427.875 0.070 428.365 ;
    RECT 0 428.435 0.070 428.925 ;
    RECT 0 428.995 0.070 429.485 ;
    RECT 0 429.555 0.070 430.045 ;
    RECT 0 430.115 0.070 430.605 ;
    RECT 0 430.675 0.070 431.165 ;
    RECT 0 431.235 0.070 431.725 ;
    RECT 0 431.795 0.070 432.285 ;
    RECT 0 432.355 0.070 432.845 ;
    RECT 0 432.915 0.070 433.405 ;
    RECT 0 433.475 0.070 433.965 ;
    RECT 0 434.035 0.070 434.525 ;
    RECT 0 434.595 0.070 435.085 ;
    RECT 0 435.155 0.070 435.645 ;
    RECT 0 435.715 0.070 436.205 ;
    RECT 0 436.275 0.070 436.765 ;
    RECT 0 436.835 0.070 437.325 ;
    RECT 0 437.395 0.070 437.885 ;
    RECT 0 437.955 0.070 438.445 ;
    RECT 0 438.515 0.070 439.005 ;
    RECT 0 439.075 0.070 439.565 ;
    RECT 0 439.635 0.070 440.125 ;
    RECT 0 440.195 0.070 440.685 ;
    RECT 0 440.755 0.070 441.245 ;
    RECT 0 441.315 0.070 441.805 ;
    RECT 0 441.875 0.070 442.365 ;
    RECT 0 442.435 0.070 442.925 ;
    RECT 0 442.995 0.070 443.485 ;
    RECT 0 443.555 0.070 444.045 ;
    RECT 0 444.115 0.070 444.605 ;
    RECT 0 444.675 0.070 445.165 ;
    RECT 0 445.235 0.070 445.725 ;
    RECT 0 445.795 0.070 446.285 ;
    RECT 0 446.355 0.070 446.845 ;
    RECT 0 446.915 0.070 447.405 ;
    RECT 0 447.475 0.070 447.965 ;
    RECT 0 448.035 0.070 448.525 ;
    RECT 0 448.595 0.070 449.085 ;
    RECT 0 449.155 0.070 449.645 ;
    RECT 0 449.715 0.070 450.205 ;
    RECT 0 450.275 0.070 450.765 ;
    RECT 0 450.835 0.070 451.325 ;
    RECT 0 451.395 0.070 451.885 ;
    RECT 0 451.955 0.070 452.445 ;
    RECT 0 452.515 0.070 453.005 ;
    RECT 0 453.075 0.070 453.565 ;
    RECT 0 453.635 0.070 454.125 ;
    RECT 0 454.195 0.070 454.685 ;
    RECT 0 454.755 0.070 455.245 ;
    RECT 0 455.315 0.070 455.805 ;
    RECT 0 455.875 0.070 456.365 ;
    RECT 0 456.435 0.070 456.925 ;
    RECT 0 456.995 0.070 457.485 ;
    RECT 0 457.555 0.070 458.045 ;
    RECT 0 458.115 0.070 458.605 ;
    RECT 0 458.675 0.070 459.165 ;
    RECT 0 459.235 0.070 459.725 ;
    RECT 0 459.795 0.070 460.285 ;
    RECT 0 460.355 0.070 460.845 ;
    RECT 0 460.915 0.070 461.405 ;
    RECT 0 461.475 0.070 461.965 ;
    RECT 0 462.035 0.070 462.525 ;
    RECT 0 462.595 0.070 463.085 ;
    RECT 0 463.155 0.070 463.645 ;
    RECT 0 463.715 0.070 464.205 ;
    RECT 0 464.275 0.070 464.765 ;
    RECT 0 464.835 0.070 465.325 ;
    RECT 0 465.395 0.070 465.885 ;
    RECT 0 465.955 0.070 466.445 ;
    RECT 0 466.515 0.070 467.005 ;
    RECT 0 467.075 0.070 467.565 ;
    RECT 0 467.635 0.070 468.125 ;
    RECT 0 468.195 0.070 468.685 ;
    RECT 0 468.755 0.070 469.245 ;
    RECT 0 469.315 0.070 469.805 ;
    RECT 0 469.875 0.070 470.365 ;
    RECT 0 470.435 0.070 470.925 ;
    RECT 0 470.995 0.070 471.485 ;
    RECT 0 471.555 0.070 472.045 ;
    RECT 0 472.115 0.070 472.605 ;
    RECT 0 472.675 0.070 473.165 ;
    RECT 0 473.235 0.070 473.725 ;
    RECT 0 473.795 0.070 474.285 ;
    RECT 0 474.355 0.070 474.845 ;
    RECT 0 474.915 0.070 475.405 ;
    RECT 0 475.475 0.070 475.965 ;
    RECT 0 476.035 0.070 476.525 ;
    RECT 0 476.595 0.070 477.085 ;
    RECT 0 477.155 0.070 477.645 ;
    RECT 0 477.715 0.070 478.205 ;
    RECT 0 478.275 0.070 478.765 ;
    RECT 0 478.835 0.070 479.325 ;
    RECT 0 479.395 0.070 479.885 ;
    RECT 0 479.955 0.070 480.445 ;
    RECT 0 480.515 0.070 481.005 ;
    RECT 0 481.075 0.070 481.565 ;
    RECT 0 481.635 0.070 482.125 ;
    RECT 0 482.195 0.070 482.685 ;
    RECT 0 482.755 0.070 483.245 ;
    RECT 0 483.315 0.070 483.805 ;
    RECT 0 483.875 0.070 484.365 ;
    RECT 0 484.435 0.070 484.925 ;
    RECT 0 484.995 0.070 485.485 ;
    RECT 0 485.555 0.070 486.045 ;
    RECT 0 486.115 0.070 486.605 ;
    RECT 0 486.675 0.070 487.165 ;
    RECT 0 487.235 0.070 487.725 ;
    RECT 0 487.795 0.070 488.285 ;
    RECT 0 488.355 0.070 488.845 ;
    RECT 0 488.915 0.070 489.405 ;
    RECT 0 489.475 0.070 489.965 ;
    RECT 0 490.035 0.070 490.525 ;
    RECT 0 490.595 0.070 491.085 ;
    RECT 0 491.155 0.070 491.645 ;
    RECT 0 491.715 0.070 492.205 ;
    RECT 0 492.275 0.070 492.765 ;
    RECT 0 492.835 0.070 493.325 ;
    RECT 0 493.395 0.070 493.885 ;
    RECT 0 493.955 0.070 494.445 ;
    RECT 0 494.515 0.070 495.005 ;
    RECT 0 495.075 0.070 495.565 ;
    RECT 0 495.635 0.070 496.125 ;
    RECT 0 496.195 0.070 496.685 ;
    RECT 0 496.755 0.070 497.245 ;
    RECT 0 497.315 0.070 497.805 ;
    RECT 0 497.875 0.070 498.365 ;
    RECT 0 498.435 0.070 498.925 ;
    RECT 0 498.995 0.070 499.485 ;
    RECT 0 499.555 0.070 500.045 ;
    RECT 0 500.115 0.070 500.605 ;
    RECT 0 500.675 0.070 501.165 ;
    RECT 0 501.235 0.070 501.725 ;
    RECT 0 501.795 0.070 502.285 ;
    RECT 0 502.355 0.070 502.845 ;
    RECT 0 502.915 0.070 503.405 ;
    RECT 0 503.475 0.070 503.965 ;
    RECT 0 504.035 0.070 504.525 ;
    RECT 0 504.595 0.070 505.085 ;
    RECT 0 505.155 0.070 505.645 ;
    RECT 0 505.715 0.070 506.205 ;
    RECT 0 506.275 0.070 506.765 ;
    RECT 0 506.835 0.070 507.325 ;
    RECT 0 507.395 0.070 507.885 ;
    RECT 0 507.955 0.070 508.445 ;
    RECT 0 508.515 0.070 509.005 ;
    RECT 0 509.075 0.070 509.565 ;
    RECT 0 509.635 0.070 510.125 ;
    RECT 0 510.195 0.070 510.685 ;
    RECT 0 510.755 0.070 511.245 ;
    RECT 0 511.315 0.070 511.805 ;
    RECT 0 511.875 0.070 512.365 ;
    RECT 0 512.435 0.070 512.925 ;
    RECT 0 512.995 0.070 513.485 ;
    RECT 0 513.555 0.070 514.045 ;
    RECT 0 514.115 0.070 514.605 ;
    RECT 0 514.675 0.070 515.165 ;
    RECT 0 515.235 0.070 515.725 ;
    RECT 0 515.795 0.070 516.285 ;
    RECT 0 516.355 0.070 516.845 ;
    RECT 0 516.915 0.070 517.405 ;
    RECT 0 517.475 0.070 517.965 ;
    RECT 0 518.035 0.070 518.525 ;
    RECT 0 518.595 0.070 519.085 ;
    RECT 0 519.155 0.070 519.645 ;
    RECT 0 519.715 0.070 520.205 ;
    RECT 0 520.275 0.070 520.765 ;
    RECT 0 520.835 0.070 521.325 ;
    RECT 0 521.395 0.070 521.885 ;
    RECT 0 521.955 0.070 522.445 ;
    RECT 0 522.515 0.070 523.005 ;
    RECT 0 523.075 0.070 523.565 ;
    RECT 0 523.635 0.070 524.125 ;
    RECT 0 524.195 0.070 524.685 ;
    RECT 0 524.755 0.070 525.245 ;
    RECT 0 525.315 0.070 525.805 ;
    RECT 0 525.875 0.070 526.365 ;
    RECT 0 526.435 0.070 526.925 ;
    RECT 0 526.995 0.070 527.485 ;
    RECT 0 527.555 0.070 528.045 ;
    RECT 0 528.115 0.070 528.605 ;
    RECT 0 528.675 0.070 529.165 ;
    RECT 0 529.235 0.070 529.725 ;
    RECT 0 529.795 0.070 530.285 ;
    RECT 0 530.355 0.070 530.845 ;
    RECT 0 530.915 0.070 531.405 ;
    RECT 0 531.475 0.070 531.965 ;
    RECT 0 532.035 0.070 532.525 ;
    RECT 0 532.595 0.070 533.085 ;
    RECT 0 533.155 0.070 533.645 ;
    RECT 0 533.715 0.070 534.205 ;
    RECT 0 534.275 0.070 534.765 ;
    RECT 0 534.835 0.070 535.325 ;
    RECT 0 535.395 0.070 535.885 ;
    RECT 0 535.955 0.070 536.445 ;
    RECT 0 536.515 0.070 537.005 ;
    RECT 0 537.075 0.070 537.565 ;
    RECT 0 537.635 0.070 538.125 ;
    RECT 0 538.195 0.070 538.685 ;
    RECT 0 538.755 0.070 539.245 ;
    RECT 0 539.315 0.070 539.805 ;
    RECT 0 539.875 0.070 540.365 ;
    RECT 0 540.435 0.070 540.925 ;
    RECT 0 540.995 0.070 541.485 ;
    RECT 0 541.555 0.070 542.045 ;
    RECT 0 542.115 0.070 542.605 ;
    RECT 0 542.675 0.070 543.165 ;
    RECT 0 543.235 0.070 543.725 ;
    RECT 0 543.795 0.070 544.285 ;
    RECT 0 544.355 0.070 544.845 ;
    RECT 0 544.915 0.070 545.405 ;
    RECT 0 545.475 0.070 545.965 ;
    RECT 0 546.035 0.070 546.525 ;
    RECT 0 546.595 0.070 547.085 ;
    RECT 0 547.155 0.070 547.645 ;
    RECT 0 547.715 0.070 548.205 ;
    RECT 0 548.275 0.070 548.765 ;
    RECT 0 548.835 0.070 549.325 ;
    RECT 0 549.395 0.070 549.885 ;
    RECT 0 549.955 0.070 550.445 ;
    RECT 0 550.515 0.070 551.005 ;
    RECT 0 551.075 0.070 551.565 ;
    RECT 0 551.635 0.070 552.125 ;
    RECT 0 552.195 0.070 552.685 ;
    RECT 0 552.755 0.070 553.245 ;
    RECT 0 553.315 0.070 553.805 ;
    RECT 0 553.875 0.070 554.365 ;
    RECT 0 554.435 0.070 554.925 ;
    RECT 0 554.995 0.070 555.485 ;
    RECT 0 555.555 0.070 556.045 ;
    RECT 0 556.115 0.070 556.605 ;
    RECT 0 556.675 0.070 557.165 ;
    RECT 0 557.235 0.070 557.725 ;
    RECT 0 557.795 0.070 558.285 ;
    RECT 0 558.355 0.070 558.845 ;
    RECT 0 558.915 0.070 559.405 ;
    RECT 0 559.475 0.070 559.965 ;
    RECT 0 560.035 0.070 560.525 ;
    RECT 0 560.595 0.070 561.085 ;
    RECT 0 561.155 0.070 561.645 ;
    RECT 0 561.715 0.070 562.205 ;
    RECT 0 562.275 0.070 562.765 ;
    RECT 0 562.835 0.070 563.325 ;
    RECT 0 563.395 0.070 563.885 ;
    RECT 0 563.955 0.070 564.445 ;
    RECT 0 564.515 0.070 565.005 ;
    RECT 0 565.075 0.070 565.565 ;
    RECT 0 565.635 0.070 566.125 ;
    RECT 0 566.195 0.070 566.685 ;
    RECT 0 566.755 0.070 567.245 ;
    RECT 0 567.315 0.070 567.805 ;
    RECT 0 567.875 0.070 568.365 ;
    RECT 0 568.435 0.070 568.925 ;
    RECT 0 568.995 0.070 569.485 ;
    RECT 0 569.555 0.070 570.045 ;
    RECT 0 570.115 0.070 570.605 ;
    RECT 0 570.675 0.070 571.165 ;
    RECT 0 571.235 0.070 571.725 ;
    RECT 0 571.795 0.070 572.285 ;
    RECT 0 572.355 0.070 572.845 ;
    RECT 0 572.915 0.070 573.405 ;
    RECT 0 573.475 0.070 573.965 ;
    RECT 0 574.035 0.070 574.525 ;
    RECT 0 574.595 0.070 575.085 ;
    RECT 0 575.155 0.070 575.645 ;
    RECT 0 575.715 0.070 576.205 ;
    RECT 0 576.275 0.070 576.765 ;
    RECT 0 576.835 0.070 577.325 ;
    RECT 0 577.395 0.070 577.885 ;
    RECT 0 577.955 0.070 578.445 ;
    RECT 0 578.515 0.070 579.005 ;
    RECT 0 579.075 0.070 579.565 ;
    RECT 0 579.635 0.070 580.125 ;
    RECT 0 580.195 0.070 580.685 ;
    RECT 0 580.755 0.070 581.245 ;
    RECT 0 581.315 0.070 581.805 ;
    RECT 0 581.875 0.070 582.365 ;
    RECT 0 582.435 0.070 582.925 ;
    RECT 0 582.995 0.070 583.485 ;
    RECT 0 583.555 0.070 584.045 ;
    RECT 0 584.115 0.070 584.605 ;
    RECT 0 584.675 0.070 585.165 ;
    RECT 0 585.235 0.070 585.725 ;
    RECT 0 585.795 0.070 586.285 ;
    RECT 0 586.355 0.070 586.845 ;
    RECT 0 586.915 0.070 587.405 ;
    RECT 0 587.475 0.070 587.965 ;
    RECT 0 588.035 0.070 588.525 ;
    RECT 0 588.595 0.070 589.085 ;
    RECT 0 589.155 0.070 589.645 ;
    RECT 0 589.715 0.070 590.205 ;
    RECT 0 590.275 0.070 590.765 ;
    RECT 0 590.835 0.070 591.325 ;
    RECT 0 591.395 0.070 591.885 ;
    RECT 0 591.955 0.070 592.445 ;
    RECT 0 592.515 0.070 593.005 ;
    RECT 0 593.075 0.070 593.565 ;
    RECT 0 593.635 0.070 594.125 ;
    RECT 0 594.195 0.070 594.685 ;
    RECT 0 594.755 0.070 595.245 ;
    RECT 0 595.315 0.070 595.805 ;
    RECT 0 595.875 0.070 596.365 ;
    RECT 0 596.435 0.070 596.925 ;
    RECT 0 596.995 0.070 597.485 ;
    RECT 0 597.555 0.070 598.045 ;
    RECT 0 598.115 0.070 598.605 ;
    RECT 0 598.675 0.070 599.165 ;
    RECT 0 599.235 0.070 599.725 ;
    RECT 0 599.795 0.070 600.285 ;
    RECT 0 600.355 0.070 600.845 ;
    RECT 0 600.915 0.070 601.405 ;
    RECT 0 601.475 0.070 629.125 ;
    RECT 0 629.195 0.070 629.685 ;
    RECT 0 629.755 0.070 630.245 ;
    RECT 0 630.315 0.070 630.805 ;
    RECT 0 630.875 0.070 631.365 ;
    RECT 0 631.435 0.070 631.925 ;
    RECT 0 631.995 0.070 632.485 ;
    RECT 0 632.555 0.070 633.045 ;
    RECT 0 633.115 0.070 633.605 ;
    RECT 0 633.675 0.070 634.165 ;
    RECT 0 634.235 0.070 634.725 ;
    RECT 0 634.795 0.070 635.285 ;
    RECT 0 635.355 0.070 635.845 ;
    RECT 0 635.915 0.070 636.405 ;
    RECT 0 636.475 0.070 636.965 ;
    RECT 0 637.035 0.070 637.525 ;
    RECT 0 637.595 0.070 638.085 ;
    RECT 0 638.155 0.070 638.645 ;
    RECT 0 638.715 0.070 639.205 ;
    RECT 0 639.275 0.070 639.765 ;
    RECT 0 639.835 0.070 640.325 ;
    RECT 0 640.395 0.070 640.885 ;
    RECT 0 640.955 0.070 641.445 ;
    RECT 0 641.515 0.070 642.005 ;
    RECT 0 642.075 0.070 642.565 ;
    RECT 0 642.635 0.070 643.125 ;
    RECT 0 643.195 0.070 643.685 ;
    RECT 0 643.755 0.070 644.245 ;
    RECT 0 644.315 0.070 644.805 ;
    RECT 0 644.875 0.070 645.365 ;
    RECT 0 645.435 0.070 645.925 ;
    RECT 0 645.995 0.070 646.485 ;
    RECT 0 646.555 0.070 647.045 ;
    RECT 0 647.115 0.070 647.605 ;
    RECT 0 647.675 0.070 648.165 ;
    RECT 0 648.235 0.070 648.725 ;
    RECT 0 648.795 0.070 649.285 ;
    RECT 0 649.355 0.070 649.845 ;
    RECT 0 649.915 0.070 650.405 ;
    RECT 0 650.475 0.070 650.965 ;
    RECT 0 651.035 0.070 651.525 ;
    RECT 0 651.595 0.070 652.085 ;
    RECT 0 652.155 0.070 652.645 ;
    RECT 0 652.715 0.070 653.205 ;
    RECT 0 653.275 0.070 653.765 ;
    RECT 0 653.835 0.070 654.325 ;
    RECT 0 654.395 0.070 654.885 ;
    RECT 0 654.955 0.070 655.445 ;
    RECT 0 655.515 0.070 656.005 ;
    RECT 0 656.075 0.070 656.565 ;
    RECT 0 656.635 0.070 657.125 ;
    RECT 0 657.195 0.070 657.685 ;
    RECT 0 657.755 0.070 658.245 ;
    RECT 0 658.315 0.070 658.805 ;
    RECT 0 658.875 0.070 659.365 ;
    RECT 0 659.435 0.070 659.925 ;
    RECT 0 659.995 0.070 660.485 ;
    RECT 0 660.555 0.070 661.045 ;
    RECT 0 661.115 0.070 661.605 ;
    RECT 0 661.675 0.070 662.165 ;
    RECT 0 662.235 0.070 662.725 ;
    RECT 0 662.795 0.070 663.285 ;
    RECT 0 663.355 0.070 663.845 ;
    RECT 0 663.915 0.070 664.405 ;
    RECT 0 664.475 0.070 664.965 ;
    RECT 0 665.035 0.070 665.525 ;
    RECT 0 665.595 0.070 666.085 ;
    RECT 0 666.155 0.070 666.645 ;
    RECT 0 666.715 0.070 667.205 ;
    RECT 0 667.275 0.070 667.765 ;
    RECT 0 667.835 0.070 668.325 ;
    RECT 0 668.395 0.070 668.885 ;
    RECT 0 668.955 0.070 669.445 ;
    RECT 0 669.515 0.070 670.005 ;
    RECT 0 670.075 0.070 670.565 ;
    RECT 0 670.635 0.070 671.125 ;
    RECT 0 671.195 0.070 671.685 ;
    RECT 0 671.755 0.070 672.245 ;
    RECT 0 672.315 0.070 672.805 ;
    RECT 0 672.875 0.070 673.365 ;
    RECT 0 673.435 0.070 673.925 ;
    RECT 0 673.995 0.070 674.485 ;
    RECT 0 674.555 0.070 675.045 ;
    RECT 0 675.115 0.070 675.605 ;
    RECT 0 675.675 0.070 676.165 ;
    RECT 0 676.235 0.070 676.725 ;
    RECT 0 676.795 0.070 677.285 ;
    RECT 0 677.355 0.070 677.845 ;
    RECT 0 677.915 0.070 678.405 ;
    RECT 0 678.475 0.070 678.965 ;
    RECT 0 679.035 0.070 679.525 ;
    RECT 0 679.595 0.070 680.085 ;
    RECT 0 680.155 0.070 680.645 ;
    RECT 0 680.715 0.070 681.205 ;
    RECT 0 681.275 0.070 681.765 ;
    RECT 0 681.835 0.070 682.325 ;
    RECT 0 682.395 0.070 682.885 ;
    RECT 0 682.955 0.070 683.445 ;
    RECT 0 683.515 0.070 684.005 ;
    RECT 0 684.075 0.070 684.565 ;
    RECT 0 684.635 0.070 685.125 ;
    RECT 0 685.195 0.070 685.685 ;
    RECT 0 685.755 0.070 686.245 ;
    RECT 0 686.315 0.070 686.805 ;
    RECT 0 686.875 0.070 687.365 ;
    RECT 0 687.435 0.070 687.925 ;
    RECT 0 687.995 0.070 688.485 ;
    RECT 0 688.555 0.070 689.045 ;
    RECT 0 689.115 0.070 689.605 ;
    RECT 0 689.675 0.070 690.165 ;
    RECT 0 690.235 0.070 690.725 ;
    RECT 0 690.795 0.070 691.285 ;
    RECT 0 691.355 0.070 691.845 ;
    RECT 0 691.915 0.070 692.405 ;
    RECT 0 692.475 0.070 692.965 ;
    RECT 0 693.035 0.070 693.525 ;
    RECT 0 693.595 0.070 694.085 ;
    RECT 0 694.155 0.070 694.645 ;
    RECT 0 694.715 0.070 695.205 ;
    RECT 0 695.275 0.070 695.765 ;
    RECT 0 695.835 0.070 696.325 ;
    RECT 0 696.395 0.070 696.885 ;
    RECT 0 696.955 0.070 697.445 ;
    RECT 0 697.515 0.070 698.005 ;
    RECT 0 698.075 0.070 698.565 ;
    RECT 0 698.635 0.070 699.125 ;
    RECT 0 699.195 0.070 699.685 ;
    RECT 0 699.755 0.070 700.245 ;
    RECT 0 700.315 0.070 700.805 ;
    RECT 0 700.875 0.070 701.365 ;
    RECT 0 701.435 0.070 701.925 ;
    RECT 0 701.995 0.070 702.485 ;
    RECT 0 702.555 0.070 703.045 ;
    RECT 0 703.115 0.070 703.605 ;
    RECT 0 703.675 0.070 704.165 ;
    RECT 0 704.235 0.070 704.725 ;
    RECT 0 704.795 0.070 705.285 ;
    RECT 0 705.355 0.070 705.845 ;
    RECT 0 705.915 0.070 706.405 ;
    RECT 0 706.475 0.070 706.965 ;
    RECT 0 707.035 0.070 707.525 ;
    RECT 0 707.595 0.070 708.085 ;
    RECT 0 708.155 0.070 708.645 ;
    RECT 0 708.715 0.070 709.205 ;
    RECT 0 709.275 0.070 709.765 ;
    RECT 0 709.835 0.070 710.325 ;
    RECT 0 710.395 0.070 710.885 ;
    RECT 0 710.955 0.070 711.445 ;
    RECT 0 711.515 0.070 712.005 ;
    RECT 0 712.075 0.070 712.565 ;
    RECT 0 712.635 0.070 713.125 ;
    RECT 0 713.195 0.070 713.685 ;
    RECT 0 713.755 0.070 714.245 ;
    RECT 0 714.315 0.070 714.805 ;
    RECT 0 714.875 0.070 715.365 ;
    RECT 0 715.435 0.070 715.925 ;
    RECT 0 715.995 0.070 716.485 ;
    RECT 0 716.555 0.070 717.045 ;
    RECT 0 717.115 0.070 717.605 ;
    RECT 0 717.675 0.070 718.165 ;
    RECT 0 718.235 0.070 718.725 ;
    RECT 0 718.795 0.070 719.285 ;
    RECT 0 719.355 0.070 719.845 ;
    RECT 0 719.915 0.070 720.405 ;
    RECT 0 720.475 0.070 720.965 ;
    RECT 0 721.035 0.070 721.525 ;
    RECT 0 721.595 0.070 722.085 ;
    RECT 0 722.155 0.070 722.645 ;
    RECT 0 722.715 0.070 723.205 ;
    RECT 0 723.275 0.070 723.765 ;
    RECT 0 723.835 0.070 724.325 ;
    RECT 0 724.395 0.070 724.885 ;
    RECT 0 724.955 0.070 725.445 ;
    RECT 0 725.515 0.070 726.005 ;
    RECT 0 726.075 0.070 726.565 ;
    RECT 0 726.635 0.070 727.125 ;
    RECT 0 727.195 0.070 727.685 ;
    RECT 0 727.755 0.070 728.245 ;
    RECT 0 728.315 0.070 728.805 ;
    RECT 0 728.875 0.070 729.365 ;
    RECT 0 729.435 0.070 729.925 ;
    RECT 0 729.995 0.070 730.485 ;
    RECT 0 730.555 0.070 731.045 ;
    RECT 0 731.115 0.070 731.605 ;
    RECT 0 731.675 0.070 732.165 ;
    RECT 0 732.235 0.070 732.725 ;
    RECT 0 732.795 0.070 733.285 ;
    RECT 0 733.355 0.070 733.845 ;
    RECT 0 733.915 0.070 734.405 ;
    RECT 0 734.475 0.070 734.965 ;
    RECT 0 735.035 0.070 735.525 ;
    RECT 0 735.595 0.070 736.085 ;
    RECT 0 736.155 0.070 736.645 ;
    RECT 0 736.715 0.070 737.205 ;
    RECT 0 737.275 0.070 737.765 ;
    RECT 0 737.835 0.070 738.325 ;
    RECT 0 738.395 0.070 738.885 ;
    RECT 0 738.955 0.070 739.445 ;
    RECT 0 739.515 0.070 740.005 ;
    RECT 0 740.075 0.070 740.565 ;
    RECT 0 740.635 0.070 741.125 ;
    RECT 0 741.195 0.070 741.685 ;
    RECT 0 741.755 0.070 742.245 ;
    RECT 0 742.315 0.070 742.805 ;
    RECT 0 742.875 0.070 743.365 ;
    RECT 0 743.435 0.070 743.925 ;
    RECT 0 743.995 0.070 744.485 ;
    RECT 0 744.555 0.070 745.045 ;
    RECT 0 745.115 0.070 745.605 ;
    RECT 0 745.675 0.070 746.165 ;
    RECT 0 746.235 0.070 746.725 ;
    RECT 0 746.795 0.070 747.285 ;
    RECT 0 747.355 0.070 747.845 ;
    RECT 0 747.915 0.070 748.405 ;
    RECT 0 748.475 0.070 748.965 ;
    RECT 0 749.035 0.070 749.525 ;
    RECT 0 749.595 0.070 750.085 ;
    RECT 0 750.155 0.070 750.645 ;
    RECT 0 750.715 0.070 751.205 ;
    RECT 0 751.275 0.070 751.765 ;
    RECT 0 751.835 0.070 752.325 ;
    RECT 0 752.395 0.070 752.885 ;
    RECT 0 752.955 0.070 753.445 ;
    RECT 0 753.515 0.070 754.005 ;
    RECT 0 754.075 0.070 754.565 ;
    RECT 0 754.635 0.070 755.125 ;
    RECT 0 755.195 0.070 755.685 ;
    RECT 0 755.755 0.070 756.245 ;
    RECT 0 756.315 0.070 756.805 ;
    RECT 0 756.875 0.070 757.365 ;
    RECT 0 757.435 0.070 757.925 ;
    RECT 0 757.995 0.070 758.485 ;
    RECT 0 758.555 0.070 759.045 ;
    RECT 0 759.115 0.070 759.605 ;
    RECT 0 759.675 0.070 760.165 ;
    RECT 0 760.235 0.070 760.725 ;
    RECT 0 760.795 0.070 761.285 ;
    RECT 0 761.355 0.070 761.845 ;
    RECT 0 761.915 0.070 762.405 ;
    RECT 0 762.475 0.070 762.965 ;
    RECT 0 763.035 0.070 763.525 ;
    RECT 0 763.595 0.070 764.085 ;
    RECT 0 764.155 0.070 764.645 ;
    RECT 0 764.715 0.070 765.205 ;
    RECT 0 765.275 0.070 765.765 ;
    RECT 0 765.835 0.070 766.325 ;
    RECT 0 766.395 0.070 766.885 ;
    RECT 0 766.955 0.070 767.445 ;
    RECT 0 767.515 0.070 768.005 ;
    RECT 0 768.075 0.070 768.565 ;
    RECT 0 768.635 0.070 769.125 ;
    RECT 0 769.195 0.070 769.685 ;
    RECT 0 769.755 0.070 770.245 ;
    RECT 0 770.315 0.070 770.805 ;
    RECT 0 770.875 0.070 771.365 ;
    RECT 0 771.435 0.070 771.925 ;
    RECT 0 771.995 0.070 772.485 ;
    RECT 0 772.555 0.070 773.045 ;
    RECT 0 773.115 0.070 773.605 ;
    RECT 0 773.675 0.070 774.165 ;
    RECT 0 774.235 0.070 774.725 ;
    RECT 0 774.795 0.070 775.285 ;
    RECT 0 775.355 0.070 775.845 ;
    RECT 0 775.915 0.070 776.405 ;
    RECT 0 776.475 0.070 776.965 ;
    RECT 0 777.035 0.070 777.525 ;
    RECT 0 777.595 0.070 778.085 ;
    RECT 0 778.155 0.070 778.645 ;
    RECT 0 778.715 0.070 779.205 ;
    RECT 0 779.275 0.070 779.765 ;
    RECT 0 779.835 0.070 780.325 ;
    RECT 0 780.395 0.070 780.885 ;
    RECT 0 780.955 0.070 781.445 ;
    RECT 0 781.515 0.070 782.005 ;
    RECT 0 782.075 0.070 782.565 ;
    RECT 0 782.635 0.070 783.125 ;
    RECT 0 783.195 0.070 783.685 ;
    RECT 0 783.755 0.070 784.245 ;
    RECT 0 784.315 0.070 784.805 ;
    RECT 0 784.875 0.070 785.365 ;
    RECT 0 785.435 0.070 785.925 ;
    RECT 0 785.995 0.070 786.485 ;
    RECT 0 786.555 0.070 787.045 ;
    RECT 0 787.115 0.070 787.605 ;
    RECT 0 787.675 0.070 788.165 ;
    RECT 0 788.235 0.070 788.725 ;
    RECT 0 788.795 0.070 789.285 ;
    RECT 0 789.355 0.070 789.845 ;
    RECT 0 789.915 0.070 790.405 ;
    RECT 0 790.475 0.070 790.965 ;
    RECT 0 791.035 0.070 791.525 ;
    RECT 0 791.595 0.070 792.085 ;
    RECT 0 792.155 0.070 792.645 ;
    RECT 0 792.715 0.070 793.205 ;
    RECT 0 793.275 0.070 793.765 ;
    RECT 0 793.835 0.070 794.325 ;
    RECT 0 794.395 0.070 794.885 ;
    RECT 0 794.955 0.070 795.445 ;
    RECT 0 795.515 0.070 796.005 ;
    RECT 0 796.075 0.070 796.565 ;
    RECT 0 796.635 0.070 797.125 ;
    RECT 0 797.195 0.070 797.685 ;
    RECT 0 797.755 0.070 798.245 ;
    RECT 0 798.315 0.070 798.805 ;
    RECT 0 798.875 0.070 799.365 ;
    RECT 0 799.435 0.070 799.925 ;
    RECT 0 799.995 0.070 800.485 ;
    RECT 0 800.555 0.070 801.045 ;
    RECT 0 801.115 0.070 801.605 ;
    RECT 0 801.675 0.070 802.165 ;
    RECT 0 802.235 0.070 802.725 ;
    RECT 0 802.795 0.070 803.285 ;
    RECT 0 803.355 0.070 803.845 ;
    RECT 0 803.915 0.070 804.405 ;
    RECT 0 804.475 0.070 804.965 ;
    RECT 0 805.035 0.070 805.525 ;
    RECT 0 805.595 0.070 806.085 ;
    RECT 0 806.155 0.070 806.645 ;
    RECT 0 806.715 0.070 807.205 ;
    RECT 0 807.275 0.070 807.765 ;
    RECT 0 807.835 0.070 808.325 ;
    RECT 0 808.395 0.070 808.885 ;
    RECT 0 808.955 0.070 809.445 ;
    RECT 0 809.515 0.070 810.005 ;
    RECT 0 810.075 0.070 810.565 ;
    RECT 0 810.635 0.070 811.125 ;
    RECT 0 811.195 0.070 811.685 ;
    RECT 0 811.755 0.070 812.245 ;
    RECT 0 812.315 0.070 812.805 ;
    RECT 0 812.875 0.070 813.365 ;
    RECT 0 813.435 0.070 813.925 ;
    RECT 0 813.995 0.070 814.485 ;
    RECT 0 814.555 0.070 815.045 ;
    RECT 0 815.115 0.070 815.605 ;
    RECT 0 815.675 0.070 816.165 ;
    RECT 0 816.235 0.070 816.725 ;
    RECT 0 816.795 0.070 817.285 ;
    RECT 0 817.355 0.070 817.845 ;
    RECT 0 817.915 0.070 818.405 ;
    RECT 0 818.475 0.070 818.965 ;
    RECT 0 819.035 0.070 819.525 ;
    RECT 0 819.595 0.070 820.085 ;
    RECT 0 820.155 0.070 820.645 ;
    RECT 0 820.715 0.070 821.205 ;
    RECT 0 821.275 0.070 821.765 ;
    RECT 0 821.835 0.070 822.325 ;
    RECT 0 822.395 0.070 822.885 ;
    RECT 0 822.955 0.070 823.445 ;
    RECT 0 823.515 0.070 824.005 ;
    RECT 0 824.075 0.070 824.565 ;
    RECT 0 824.635 0.070 825.125 ;
    RECT 0 825.195 0.070 825.685 ;
    RECT 0 825.755 0.070 826.245 ;
    RECT 0 826.315 0.070 826.805 ;
    RECT 0 826.875 0.070 827.365 ;
    RECT 0 827.435 0.070 827.925 ;
    RECT 0 827.995 0.070 828.485 ;
    RECT 0 828.555 0.070 829.045 ;
    RECT 0 829.115 0.070 829.605 ;
    RECT 0 829.675 0.070 830.165 ;
    RECT 0 830.235 0.070 830.725 ;
    RECT 0 830.795 0.070 831.285 ;
    RECT 0 831.355 0.070 831.845 ;
    RECT 0 831.915 0.070 832.405 ;
    RECT 0 832.475 0.070 832.965 ;
    RECT 0 833.035 0.070 833.525 ;
    RECT 0 833.595 0.070 834.085 ;
    RECT 0 834.155 0.070 834.645 ;
    RECT 0 834.715 0.070 835.205 ;
    RECT 0 835.275 0.070 835.765 ;
    RECT 0 835.835 0.070 836.325 ;
    RECT 0 836.395 0.070 836.885 ;
    RECT 0 836.955 0.070 837.445 ;
    RECT 0 837.515 0.070 838.005 ;
    RECT 0 838.075 0.070 838.565 ;
    RECT 0 838.635 0.070 839.125 ;
    RECT 0 839.195 0.070 839.685 ;
    RECT 0 839.755 0.070 840.245 ;
    RECT 0 840.315 0.070 840.805 ;
    RECT 0 840.875 0.070 841.365 ;
    RECT 0 841.435 0.070 841.925 ;
    RECT 0 841.995 0.070 842.485 ;
    RECT 0 842.555 0.070 843.045 ;
    RECT 0 843.115 0.070 843.605 ;
    RECT 0 843.675 0.070 844.165 ;
    RECT 0 844.235 0.070 844.725 ;
    RECT 0 844.795 0.070 845.285 ;
    RECT 0 845.355 0.070 845.845 ;
    RECT 0 845.915 0.070 846.405 ;
    RECT 0 846.475 0.070 846.965 ;
    RECT 0 847.035 0.070 847.525 ;
    RECT 0 847.595 0.070 848.085 ;
    RECT 0 848.155 0.070 848.645 ;
    RECT 0 848.715 0.070 849.205 ;
    RECT 0 849.275 0.070 849.765 ;
    RECT 0 849.835 0.070 850.325 ;
    RECT 0 850.395 0.070 850.885 ;
    RECT 0 850.955 0.070 851.445 ;
    RECT 0 851.515 0.070 852.005 ;
    RECT 0 852.075 0.070 852.565 ;
    RECT 0 852.635 0.070 853.125 ;
    RECT 0 853.195 0.070 853.685 ;
    RECT 0 853.755 0.070 854.245 ;
    RECT 0 854.315 0.070 854.805 ;
    RECT 0 854.875 0.070 855.365 ;
    RECT 0 855.435 0.070 855.925 ;
    RECT 0 855.995 0.070 856.485 ;
    RECT 0 856.555 0.070 857.045 ;
    RECT 0 857.115 0.070 857.605 ;
    RECT 0 857.675 0.070 858.165 ;
    RECT 0 858.235 0.070 858.725 ;
    RECT 0 858.795 0.070 859.285 ;
    RECT 0 859.355 0.070 859.845 ;
    RECT 0 859.915 0.070 860.405 ;
    RECT 0 860.475 0.070 860.965 ;
    RECT 0 861.035 0.070 861.525 ;
    RECT 0 861.595 0.070 862.085 ;
    RECT 0 862.155 0.070 862.645 ;
    RECT 0 862.715 0.070 863.205 ;
    RECT 0 863.275 0.070 863.765 ;
    RECT 0 863.835 0.070 864.325 ;
    RECT 0 864.395 0.070 864.885 ;
    RECT 0 864.955 0.070 865.445 ;
    RECT 0 865.515 0.070 866.005 ;
    RECT 0 866.075 0.070 866.565 ;
    RECT 0 866.635 0.070 867.125 ;
    RECT 0 867.195 0.070 867.685 ;
    RECT 0 867.755 0.070 868.245 ;
    RECT 0 868.315 0.070 868.805 ;
    RECT 0 868.875 0.070 869.365 ;
    RECT 0 869.435 0.070 869.925 ;
    RECT 0 869.995 0.070 870.485 ;
    RECT 0 870.555 0.070 871.045 ;
    RECT 0 871.115 0.070 871.605 ;
    RECT 0 871.675 0.070 872.165 ;
    RECT 0 872.235 0.070 872.725 ;
    RECT 0 872.795 0.070 873.285 ;
    RECT 0 873.355 0.070 873.845 ;
    RECT 0 873.915 0.070 874.405 ;
    RECT 0 874.475 0.070 874.965 ;
    RECT 0 875.035 0.070 875.525 ;
    RECT 0 875.595 0.070 876.085 ;
    RECT 0 876.155 0.070 876.645 ;
    RECT 0 876.715 0.070 877.205 ;
    RECT 0 877.275 0.070 877.765 ;
    RECT 0 877.835 0.070 878.325 ;
    RECT 0 878.395 0.070 878.885 ;
    RECT 0 878.955 0.070 879.445 ;
    RECT 0 879.515 0.070 880.005 ;
    RECT 0 880.075 0.070 880.565 ;
    RECT 0 880.635 0.070 881.125 ;
    RECT 0 881.195 0.070 881.685 ;
    RECT 0 881.755 0.070 882.245 ;
    RECT 0 882.315 0.070 882.805 ;
    RECT 0 882.875 0.070 883.365 ;
    RECT 0 883.435 0.070 883.925 ;
    RECT 0 883.995 0.070 884.485 ;
    RECT 0 884.555 0.070 885.045 ;
    RECT 0 885.115 0.070 885.605 ;
    RECT 0 885.675 0.070 886.165 ;
    RECT 0 886.235 0.070 886.725 ;
    RECT 0 886.795 0.070 887.285 ;
    RECT 0 887.355 0.070 887.845 ;
    RECT 0 887.915 0.070 888.405 ;
    RECT 0 888.475 0.070 888.965 ;
    RECT 0 889.035 0.070 889.525 ;
    RECT 0 889.595 0.070 890.085 ;
    RECT 0 890.155 0.070 890.645 ;
    RECT 0 890.715 0.070 891.205 ;
    RECT 0 891.275 0.070 891.765 ;
    RECT 0 891.835 0.070 892.325 ;
    RECT 0 892.395 0.070 892.885 ;
    RECT 0 892.955 0.070 893.445 ;
    RECT 0 893.515 0.070 894.005 ;
    RECT 0 894.075 0.070 894.565 ;
    RECT 0 894.635 0.070 895.125 ;
    RECT 0 895.195 0.070 895.685 ;
    RECT 0 895.755 0.070 896.245 ;
    RECT 0 896.315 0.070 896.805 ;
    RECT 0 896.875 0.070 897.365 ;
    RECT 0 897.435 0.070 897.925 ;
    RECT 0 897.995 0.070 898.485 ;
    RECT 0 898.555 0.070 899.045 ;
    RECT 0 899.115 0.070 899.605 ;
    RECT 0 899.675 0.070 900.165 ;
    RECT 0 900.235 0.070 900.725 ;
    RECT 0 900.795 0.070 901.285 ;
    RECT 0 901.355 0.070 901.845 ;
    RECT 0 901.915 0.070 902.405 ;
    RECT 0 902.475 0.070 902.965 ;
    RECT 0 903.035 0.070 903.525 ;
    RECT 0 903.595 0.070 904.085 ;
    RECT 0 904.155 0.070 904.645 ;
    RECT 0 904.715 0.070 905.205 ;
    RECT 0 905.275 0.070 905.765 ;
    RECT 0 905.835 0.070 906.325 ;
    RECT 0 906.395 0.070 906.885 ;
    RECT 0 906.955 0.070 907.445 ;
    RECT 0 907.515 0.070 908.005 ;
    RECT 0 908.075 0.070 908.565 ;
    RECT 0 908.635 0.070 909.125 ;
    RECT 0 909.195 0.070 909.685 ;
    RECT 0 909.755 0.070 910.245 ;
    RECT 0 910.315 0.070 910.805 ;
    RECT 0 910.875 0.070 911.365 ;
    RECT 0 911.435 0.070 911.925 ;
    RECT 0 911.995 0.070 912.485 ;
    RECT 0 912.555 0.070 913.045 ;
    RECT 0 913.115 0.070 913.605 ;
    RECT 0 913.675 0.070 914.165 ;
    RECT 0 914.235 0.070 914.725 ;
    RECT 0 914.795 0.070 915.285 ;
    RECT 0 915.355 0.070 943.005 ;
    RECT 0 943.075 0.070 943.565 ;
    RECT 0 943.635 0.070 944.125 ;
    RECT 0 944.195 0.070 944.685 ;
    RECT 0 944.755 0.070 945.245 ;
    RECT 0 945.315 0.070 945.805 ;
    RECT 0 945.875 0.070 946.365 ;
    RECT 0 946.435 0.070 946.925 ;
    RECT 0 946.995 0.070 947.485 ;
    RECT 0 947.555 0.070 948.045 ;
    RECT 0 948.115 0.070 975.765 ;
    RECT 0 975.835 0.070 976.325 ;
    RECT 0 976.395 0.070 976.885 ;
    RECT 0 976.955 0.070 981.400 ;
    LAYER metal4 ;
    RECT 0 0 1832.740 1.400 ;
    RECT 0 980.000 1832.740 981.400 ;
    RECT 0.000 1.400 1.260 980.000 ;
    RECT 1.540 1.400 2.380 980.000 ;
    RECT 2.660 1.400 3.500 980.000 ;
    RECT 3.780 1.400 4.620 980.000 ;
    RECT 4.900 1.400 5.740 980.000 ;
    RECT 6.020 1.400 6.860 980.000 ;
    RECT 7.140 1.400 7.980 980.000 ;
    RECT 8.260 1.400 9.100 980.000 ;
    RECT 9.380 1.400 10.220 980.000 ;
    RECT 10.500 1.400 11.340 980.000 ;
    RECT 11.620 1.400 12.460 980.000 ;
    RECT 12.740 1.400 13.580 980.000 ;
    RECT 13.860 1.400 14.700 980.000 ;
    RECT 14.980 1.400 15.820 980.000 ;
    RECT 16.100 1.400 16.940 980.000 ;
    RECT 17.220 1.400 18.060 980.000 ;
    RECT 18.340 1.400 19.180 980.000 ;
    RECT 19.460 1.400 20.300 980.000 ;
    RECT 20.580 1.400 21.420 980.000 ;
    RECT 21.700 1.400 22.540 980.000 ;
    RECT 22.820 1.400 23.660 980.000 ;
    RECT 23.940 1.400 24.780 980.000 ;
    RECT 25.060 1.400 25.900 980.000 ;
    RECT 26.180 1.400 27.020 980.000 ;
    RECT 27.300 1.400 28.140 980.000 ;
    RECT 28.420 1.400 29.260 980.000 ;
    RECT 29.540 1.400 30.380 980.000 ;
    RECT 30.660 1.400 31.500 980.000 ;
    RECT 31.780 1.400 32.620 980.000 ;
    RECT 32.900 1.400 33.740 980.000 ;
    RECT 34.020 1.400 34.860 980.000 ;
    RECT 35.140 1.400 35.980 980.000 ;
    RECT 36.260 1.400 37.100 980.000 ;
    RECT 37.380 1.400 38.220 980.000 ;
    RECT 38.500 1.400 39.340 980.000 ;
    RECT 39.620 1.400 40.460 980.000 ;
    RECT 40.740 1.400 41.580 980.000 ;
    RECT 41.860 1.400 42.700 980.000 ;
    RECT 42.980 1.400 43.820 980.000 ;
    RECT 44.100 1.400 44.940 980.000 ;
    RECT 45.220 1.400 46.060 980.000 ;
    RECT 46.340 1.400 47.180 980.000 ;
    RECT 47.460 1.400 48.300 980.000 ;
    RECT 48.580 1.400 49.420 980.000 ;
    RECT 49.700 1.400 50.540 980.000 ;
    RECT 50.820 1.400 51.660 980.000 ;
    RECT 51.940 1.400 52.780 980.000 ;
    RECT 53.060 1.400 53.900 980.000 ;
    RECT 54.180 1.400 55.020 980.000 ;
    RECT 55.300 1.400 56.140 980.000 ;
    RECT 56.420 1.400 57.260 980.000 ;
    RECT 57.540 1.400 58.380 980.000 ;
    RECT 58.660 1.400 59.500 980.000 ;
    RECT 59.780 1.400 60.620 980.000 ;
    RECT 60.900 1.400 61.740 980.000 ;
    RECT 62.020 1.400 62.860 980.000 ;
    RECT 63.140 1.400 63.980 980.000 ;
    RECT 64.260 1.400 65.100 980.000 ;
    RECT 65.380 1.400 66.220 980.000 ;
    RECT 66.500 1.400 67.340 980.000 ;
    RECT 67.620 1.400 68.460 980.000 ;
    RECT 68.740 1.400 69.580 980.000 ;
    RECT 69.860 1.400 70.700 980.000 ;
    RECT 70.980 1.400 71.820 980.000 ;
    RECT 72.100 1.400 72.940 980.000 ;
    RECT 73.220 1.400 74.060 980.000 ;
    RECT 74.340 1.400 75.180 980.000 ;
    RECT 75.460 1.400 76.300 980.000 ;
    RECT 76.580 1.400 77.420 980.000 ;
    RECT 77.700 1.400 78.540 980.000 ;
    RECT 78.820 1.400 79.660 980.000 ;
    RECT 79.940 1.400 80.780 980.000 ;
    RECT 81.060 1.400 81.900 980.000 ;
    RECT 82.180 1.400 83.020 980.000 ;
    RECT 83.300 1.400 84.140 980.000 ;
    RECT 84.420 1.400 85.260 980.000 ;
    RECT 85.540 1.400 86.380 980.000 ;
    RECT 86.660 1.400 87.500 980.000 ;
    RECT 87.780 1.400 88.620 980.000 ;
    RECT 88.900 1.400 89.740 980.000 ;
    RECT 90.020 1.400 90.860 980.000 ;
    RECT 91.140 1.400 91.980 980.000 ;
    RECT 92.260 1.400 93.100 980.000 ;
    RECT 93.380 1.400 94.220 980.000 ;
    RECT 94.500 1.400 95.340 980.000 ;
    RECT 95.620 1.400 96.460 980.000 ;
    RECT 96.740 1.400 97.580 980.000 ;
    RECT 97.860 1.400 98.700 980.000 ;
    RECT 98.980 1.400 99.820 980.000 ;
    RECT 100.100 1.400 100.940 980.000 ;
    RECT 101.220 1.400 102.060 980.000 ;
    RECT 102.340 1.400 103.180 980.000 ;
    RECT 103.460 1.400 104.300 980.000 ;
    RECT 104.580 1.400 105.420 980.000 ;
    RECT 105.700 1.400 106.540 980.000 ;
    RECT 106.820 1.400 107.660 980.000 ;
    RECT 107.940 1.400 108.780 980.000 ;
    RECT 109.060 1.400 109.900 980.000 ;
    RECT 110.180 1.400 111.020 980.000 ;
    RECT 111.300 1.400 112.140 980.000 ;
    RECT 112.420 1.400 113.260 980.000 ;
    RECT 113.540 1.400 114.380 980.000 ;
    RECT 114.660 1.400 115.500 980.000 ;
    RECT 115.780 1.400 116.620 980.000 ;
    RECT 116.900 1.400 117.740 980.000 ;
    RECT 118.020 1.400 118.860 980.000 ;
    RECT 119.140 1.400 119.980 980.000 ;
    RECT 120.260 1.400 121.100 980.000 ;
    RECT 121.380 1.400 122.220 980.000 ;
    RECT 122.500 1.400 123.340 980.000 ;
    RECT 123.620 1.400 124.460 980.000 ;
    RECT 124.740 1.400 125.580 980.000 ;
    RECT 125.860 1.400 126.700 980.000 ;
    RECT 126.980 1.400 127.820 980.000 ;
    RECT 128.100 1.400 128.940 980.000 ;
    RECT 129.220 1.400 130.060 980.000 ;
    RECT 130.340 1.400 131.180 980.000 ;
    RECT 131.460 1.400 132.300 980.000 ;
    RECT 132.580 1.400 133.420 980.000 ;
    RECT 133.700 1.400 134.540 980.000 ;
    RECT 134.820 1.400 135.660 980.000 ;
    RECT 135.940 1.400 136.780 980.000 ;
    RECT 137.060 1.400 137.900 980.000 ;
    RECT 138.180 1.400 139.020 980.000 ;
    RECT 139.300 1.400 140.140 980.000 ;
    RECT 140.420 1.400 141.260 980.000 ;
    RECT 141.540 1.400 142.380 980.000 ;
    RECT 142.660 1.400 143.500 980.000 ;
    RECT 143.780 1.400 144.620 980.000 ;
    RECT 144.900 1.400 145.740 980.000 ;
    RECT 146.020 1.400 146.860 980.000 ;
    RECT 147.140 1.400 147.980 980.000 ;
    RECT 148.260 1.400 149.100 980.000 ;
    RECT 149.380 1.400 150.220 980.000 ;
    RECT 150.500 1.400 151.340 980.000 ;
    RECT 151.620 1.400 152.460 980.000 ;
    RECT 152.740 1.400 153.580 980.000 ;
    RECT 153.860 1.400 154.700 980.000 ;
    RECT 154.980 1.400 155.820 980.000 ;
    RECT 156.100 1.400 156.940 980.000 ;
    RECT 157.220 1.400 158.060 980.000 ;
    RECT 158.340 1.400 159.180 980.000 ;
    RECT 159.460 1.400 160.300 980.000 ;
    RECT 160.580 1.400 161.420 980.000 ;
    RECT 161.700 1.400 162.540 980.000 ;
    RECT 162.820 1.400 163.660 980.000 ;
    RECT 163.940 1.400 164.780 980.000 ;
    RECT 165.060 1.400 165.900 980.000 ;
    RECT 166.180 1.400 167.020 980.000 ;
    RECT 167.300 1.400 168.140 980.000 ;
    RECT 168.420 1.400 169.260 980.000 ;
    RECT 169.540 1.400 170.380 980.000 ;
    RECT 170.660 1.400 171.500 980.000 ;
    RECT 171.780 1.400 172.620 980.000 ;
    RECT 172.900 1.400 173.740 980.000 ;
    RECT 174.020 1.400 174.860 980.000 ;
    RECT 175.140 1.400 175.980 980.000 ;
    RECT 176.260 1.400 177.100 980.000 ;
    RECT 177.380 1.400 178.220 980.000 ;
    RECT 178.500 1.400 179.340 980.000 ;
    RECT 179.620 1.400 180.460 980.000 ;
    RECT 180.740 1.400 181.580 980.000 ;
    RECT 181.860 1.400 182.700 980.000 ;
    RECT 182.980 1.400 183.820 980.000 ;
    RECT 184.100 1.400 184.940 980.000 ;
    RECT 185.220 1.400 186.060 980.000 ;
    RECT 186.340 1.400 187.180 980.000 ;
    RECT 187.460 1.400 188.300 980.000 ;
    RECT 188.580 1.400 189.420 980.000 ;
    RECT 189.700 1.400 190.540 980.000 ;
    RECT 190.820 1.400 191.660 980.000 ;
    RECT 191.940 1.400 192.780 980.000 ;
    RECT 193.060 1.400 193.900 980.000 ;
    RECT 194.180 1.400 195.020 980.000 ;
    RECT 195.300 1.400 196.140 980.000 ;
    RECT 196.420 1.400 197.260 980.000 ;
    RECT 197.540 1.400 198.380 980.000 ;
    RECT 198.660 1.400 199.500 980.000 ;
    RECT 199.780 1.400 200.620 980.000 ;
    RECT 200.900 1.400 201.740 980.000 ;
    RECT 202.020 1.400 202.860 980.000 ;
    RECT 203.140 1.400 203.980 980.000 ;
    RECT 204.260 1.400 205.100 980.000 ;
    RECT 205.380 1.400 206.220 980.000 ;
    RECT 206.500 1.400 207.340 980.000 ;
    RECT 207.620 1.400 208.460 980.000 ;
    RECT 208.740 1.400 209.580 980.000 ;
    RECT 209.860 1.400 210.700 980.000 ;
    RECT 210.980 1.400 211.820 980.000 ;
    RECT 212.100 1.400 212.940 980.000 ;
    RECT 213.220 1.400 214.060 980.000 ;
    RECT 214.340 1.400 215.180 980.000 ;
    RECT 215.460 1.400 216.300 980.000 ;
    RECT 216.580 1.400 217.420 980.000 ;
    RECT 217.700 1.400 218.540 980.000 ;
    RECT 218.820 1.400 219.660 980.000 ;
    RECT 219.940 1.400 220.780 980.000 ;
    RECT 221.060 1.400 221.900 980.000 ;
    RECT 222.180 1.400 223.020 980.000 ;
    RECT 223.300 1.400 224.140 980.000 ;
    RECT 224.420 1.400 225.260 980.000 ;
    RECT 225.540 1.400 226.380 980.000 ;
    RECT 226.660 1.400 227.500 980.000 ;
    RECT 227.780 1.400 228.620 980.000 ;
    RECT 228.900 1.400 229.740 980.000 ;
    RECT 230.020 1.400 230.860 980.000 ;
    RECT 231.140 1.400 231.980 980.000 ;
    RECT 232.260 1.400 233.100 980.000 ;
    RECT 233.380 1.400 234.220 980.000 ;
    RECT 234.500 1.400 235.340 980.000 ;
    RECT 235.620 1.400 236.460 980.000 ;
    RECT 236.740 1.400 237.580 980.000 ;
    RECT 237.860 1.400 238.700 980.000 ;
    RECT 238.980 1.400 239.820 980.000 ;
    RECT 240.100 1.400 240.940 980.000 ;
    RECT 241.220 1.400 242.060 980.000 ;
    RECT 242.340 1.400 243.180 980.000 ;
    RECT 243.460 1.400 244.300 980.000 ;
    RECT 244.580 1.400 245.420 980.000 ;
    RECT 245.700 1.400 246.540 980.000 ;
    RECT 246.820 1.400 247.660 980.000 ;
    RECT 247.940 1.400 248.780 980.000 ;
    RECT 249.060 1.400 249.900 980.000 ;
    RECT 250.180 1.400 251.020 980.000 ;
    RECT 251.300 1.400 252.140 980.000 ;
    RECT 252.420 1.400 253.260 980.000 ;
    RECT 253.540 1.400 254.380 980.000 ;
    RECT 254.660 1.400 255.500 980.000 ;
    RECT 255.780 1.400 256.620 980.000 ;
    RECT 256.900 1.400 257.740 980.000 ;
    RECT 258.020 1.400 258.860 980.000 ;
    RECT 259.140 1.400 259.980 980.000 ;
    RECT 260.260 1.400 261.100 980.000 ;
    RECT 261.380 1.400 262.220 980.000 ;
    RECT 262.500 1.400 263.340 980.000 ;
    RECT 263.620 1.400 264.460 980.000 ;
    RECT 264.740 1.400 265.580 980.000 ;
    RECT 265.860 1.400 266.700 980.000 ;
    RECT 266.980 1.400 267.820 980.000 ;
    RECT 268.100 1.400 268.940 980.000 ;
    RECT 269.220 1.400 270.060 980.000 ;
    RECT 270.340 1.400 271.180 980.000 ;
    RECT 271.460 1.400 272.300 980.000 ;
    RECT 272.580 1.400 273.420 980.000 ;
    RECT 273.700 1.400 274.540 980.000 ;
    RECT 274.820 1.400 275.660 980.000 ;
    RECT 275.940 1.400 276.780 980.000 ;
    RECT 277.060 1.400 277.900 980.000 ;
    RECT 278.180 1.400 279.020 980.000 ;
    RECT 279.300 1.400 280.140 980.000 ;
    RECT 280.420 1.400 281.260 980.000 ;
    RECT 281.540 1.400 282.380 980.000 ;
    RECT 282.660 1.400 283.500 980.000 ;
    RECT 283.780 1.400 284.620 980.000 ;
    RECT 284.900 1.400 285.740 980.000 ;
    RECT 286.020 1.400 286.860 980.000 ;
    RECT 287.140 1.400 287.980 980.000 ;
    RECT 288.260 1.400 289.100 980.000 ;
    RECT 289.380 1.400 290.220 980.000 ;
    RECT 290.500 1.400 291.340 980.000 ;
    RECT 291.620 1.400 292.460 980.000 ;
    RECT 292.740 1.400 293.580 980.000 ;
    RECT 293.860 1.400 294.700 980.000 ;
    RECT 294.980 1.400 295.820 980.000 ;
    RECT 296.100 1.400 296.940 980.000 ;
    RECT 297.220 1.400 298.060 980.000 ;
    RECT 298.340 1.400 299.180 980.000 ;
    RECT 299.460 1.400 300.300 980.000 ;
    RECT 300.580 1.400 301.420 980.000 ;
    RECT 301.700 1.400 302.540 980.000 ;
    RECT 302.820 1.400 303.660 980.000 ;
    RECT 303.940 1.400 304.780 980.000 ;
    RECT 305.060 1.400 305.900 980.000 ;
    RECT 306.180 1.400 307.020 980.000 ;
    RECT 307.300 1.400 308.140 980.000 ;
    RECT 308.420 1.400 309.260 980.000 ;
    RECT 309.540 1.400 310.380 980.000 ;
    RECT 310.660 1.400 311.500 980.000 ;
    RECT 311.780 1.400 312.620 980.000 ;
    RECT 312.900 1.400 313.740 980.000 ;
    RECT 314.020 1.400 314.860 980.000 ;
    RECT 315.140 1.400 315.980 980.000 ;
    RECT 316.260 1.400 317.100 980.000 ;
    RECT 317.380 1.400 318.220 980.000 ;
    RECT 318.500 1.400 319.340 980.000 ;
    RECT 319.620 1.400 320.460 980.000 ;
    RECT 320.740 1.400 321.580 980.000 ;
    RECT 321.860 1.400 322.700 980.000 ;
    RECT 322.980 1.400 323.820 980.000 ;
    RECT 324.100 1.400 324.940 980.000 ;
    RECT 325.220 1.400 326.060 980.000 ;
    RECT 326.340 1.400 327.180 980.000 ;
    RECT 327.460 1.400 328.300 980.000 ;
    RECT 328.580 1.400 329.420 980.000 ;
    RECT 329.700 1.400 330.540 980.000 ;
    RECT 330.820 1.400 331.660 980.000 ;
    RECT 331.940 1.400 332.780 980.000 ;
    RECT 333.060 1.400 333.900 980.000 ;
    RECT 334.180 1.400 335.020 980.000 ;
    RECT 335.300 1.400 336.140 980.000 ;
    RECT 336.420 1.400 337.260 980.000 ;
    RECT 337.540 1.400 338.380 980.000 ;
    RECT 338.660 1.400 339.500 980.000 ;
    RECT 339.780 1.400 340.620 980.000 ;
    RECT 340.900 1.400 341.740 980.000 ;
    RECT 342.020 1.400 342.860 980.000 ;
    RECT 343.140 1.400 343.980 980.000 ;
    RECT 344.260 1.400 345.100 980.000 ;
    RECT 345.380 1.400 346.220 980.000 ;
    RECT 346.500 1.400 347.340 980.000 ;
    RECT 347.620 1.400 348.460 980.000 ;
    RECT 348.740 1.400 349.580 980.000 ;
    RECT 349.860 1.400 350.700 980.000 ;
    RECT 350.980 1.400 351.820 980.000 ;
    RECT 352.100 1.400 352.940 980.000 ;
    RECT 353.220 1.400 354.060 980.000 ;
    RECT 354.340 1.400 355.180 980.000 ;
    RECT 355.460 1.400 356.300 980.000 ;
    RECT 356.580 1.400 357.420 980.000 ;
    RECT 357.700 1.400 358.540 980.000 ;
    RECT 358.820 1.400 359.660 980.000 ;
    RECT 359.940 1.400 360.780 980.000 ;
    RECT 361.060 1.400 361.900 980.000 ;
    RECT 362.180 1.400 363.020 980.000 ;
    RECT 363.300 1.400 364.140 980.000 ;
    RECT 364.420 1.400 365.260 980.000 ;
    RECT 365.540 1.400 366.380 980.000 ;
    RECT 366.660 1.400 367.500 980.000 ;
    RECT 367.780 1.400 368.620 980.000 ;
    RECT 368.900 1.400 369.740 980.000 ;
    RECT 370.020 1.400 370.860 980.000 ;
    RECT 371.140 1.400 371.980 980.000 ;
    RECT 372.260 1.400 373.100 980.000 ;
    RECT 373.380 1.400 374.220 980.000 ;
    RECT 374.500 1.400 375.340 980.000 ;
    RECT 375.620 1.400 376.460 980.000 ;
    RECT 376.740 1.400 377.580 980.000 ;
    RECT 377.860 1.400 378.700 980.000 ;
    RECT 378.980 1.400 379.820 980.000 ;
    RECT 380.100 1.400 380.940 980.000 ;
    RECT 381.220 1.400 382.060 980.000 ;
    RECT 382.340 1.400 383.180 980.000 ;
    RECT 383.460 1.400 384.300 980.000 ;
    RECT 384.580 1.400 385.420 980.000 ;
    RECT 385.700 1.400 386.540 980.000 ;
    RECT 386.820 1.400 387.660 980.000 ;
    RECT 387.940 1.400 388.780 980.000 ;
    RECT 389.060 1.400 389.900 980.000 ;
    RECT 390.180 1.400 391.020 980.000 ;
    RECT 391.300 1.400 392.140 980.000 ;
    RECT 392.420 1.400 393.260 980.000 ;
    RECT 393.540 1.400 394.380 980.000 ;
    RECT 394.660 1.400 395.500 980.000 ;
    RECT 395.780 1.400 396.620 980.000 ;
    RECT 396.900 1.400 397.740 980.000 ;
    RECT 398.020 1.400 398.860 980.000 ;
    RECT 399.140 1.400 399.980 980.000 ;
    RECT 400.260 1.400 401.100 980.000 ;
    RECT 401.380 1.400 402.220 980.000 ;
    RECT 402.500 1.400 403.340 980.000 ;
    RECT 403.620 1.400 404.460 980.000 ;
    RECT 404.740 1.400 405.580 980.000 ;
    RECT 405.860 1.400 406.700 980.000 ;
    RECT 406.980 1.400 407.820 980.000 ;
    RECT 408.100 1.400 408.940 980.000 ;
    RECT 409.220 1.400 410.060 980.000 ;
    RECT 410.340 1.400 411.180 980.000 ;
    RECT 411.460 1.400 412.300 980.000 ;
    RECT 412.580 1.400 413.420 980.000 ;
    RECT 413.700 1.400 414.540 980.000 ;
    RECT 414.820 1.400 415.660 980.000 ;
    RECT 415.940 1.400 416.780 980.000 ;
    RECT 417.060 1.400 417.900 980.000 ;
    RECT 418.180 1.400 419.020 980.000 ;
    RECT 419.300 1.400 420.140 980.000 ;
    RECT 420.420 1.400 421.260 980.000 ;
    RECT 421.540 1.400 422.380 980.000 ;
    RECT 422.660 1.400 423.500 980.000 ;
    RECT 423.780 1.400 424.620 980.000 ;
    RECT 424.900 1.400 425.740 980.000 ;
    RECT 426.020 1.400 426.860 980.000 ;
    RECT 427.140 1.400 427.980 980.000 ;
    RECT 428.260 1.400 429.100 980.000 ;
    RECT 429.380 1.400 430.220 980.000 ;
    RECT 430.500 1.400 431.340 980.000 ;
    RECT 431.620 1.400 432.460 980.000 ;
    RECT 432.740 1.400 433.580 980.000 ;
    RECT 433.860 1.400 434.700 980.000 ;
    RECT 434.980 1.400 435.820 980.000 ;
    RECT 436.100 1.400 436.940 980.000 ;
    RECT 437.220 1.400 438.060 980.000 ;
    RECT 438.340 1.400 439.180 980.000 ;
    RECT 439.460 1.400 440.300 980.000 ;
    RECT 440.580 1.400 441.420 980.000 ;
    RECT 441.700 1.400 442.540 980.000 ;
    RECT 442.820 1.400 443.660 980.000 ;
    RECT 443.940 1.400 444.780 980.000 ;
    RECT 445.060 1.400 445.900 980.000 ;
    RECT 446.180 1.400 447.020 980.000 ;
    RECT 447.300 1.400 448.140 980.000 ;
    RECT 448.420 1.400 449.260 980.000 ;
    RECT 449.540 1.400 450.380 980.000 ;
    RECT 450.660 1.400 451.500 980.000 ;
    RECT 451.780 1.400 452.620 980.000 ;
    RECT 452.900 1.400 453.740 980.000 ;
    RECT 454.020 1.400 454.860 980.000 ;
    RECT 455.140 1.400 455.980 980.000 ;
    RECT 456.260 1.400 457.100 980.000 ;
    RECT 457.380 1.400 458.220 980.000 ;
    RECT 458.500 1.400 459.340 980.000 ;
    RECT 459.620 1.400 460.460 980.000 ;
    RECT 460.740 1.400 461.580 980.000 ;
    RECT 461.860 1.400 462.700 980.000 ;
    RECT 462.980 1.400 463.820 980.000 ;
    RECT 464.100 1.400 464.940 980.000 ;
    RECT 465.220 1.400 466.060 980.000 ;
    RECT 466.340 1.400 467.180 980.000 ;
    RECT 467.460 1.400 468.300 980.000 ;
    RECT 468.580 1.400 469.420 980.000 ;
    RECT 469.700 1.400 470.540 980.000 ;
    RECT 470.820 1.400 471.660 980.000 ;
    RECT 471.940 1.400 472.780 980.000 ;
    RECT 473.060 1.400 473.900 980.000 ;
    RECT 474.180 1.400 475.020 980.000 ;
    RECT 475.300 1.400 476.140 980.000 ;
    RECT 476.420 1.400 477.260 980.000 ;
    RECT 477.540 1.400 478.380 980.000 ;
    RECT 478.660 1.400 479.500 980.000 ;
    RECT 479.780 1.400 480.620 980.000 ;
    RECT 480.900 1.400 481.740 980.000 ;
    RECT 482.020 1.400 482.860 980.000 ;
    RECT 483.140 1.400 483.980 980.000 ;
    RECT 484.260 1.400 485.100 980.000 ;
    RECT 485.380 1.400 486.220 980.000 ;
    RECT 486.500 1.400 487.340 980.000 ;
    RECT 487.620 1.400 488.460 980.000 ;
    RECT 488.740 1.400 489.580 980.000 ;
    RECT 489.860 1.400 490.700 980.000 ;
    RECT 490.980 1.400 491.820 980.000 ;
    RECT 492.100 1.400 492.940 980.000 ;
    RECT 493.220 1.400 494.060 980.000 ;
    RECT 494.340 1.400 495.180 980.000 ;
    RECT 495.460 1.400 496.300 980.000 ;
    RECT 496.580 1.400 497.420 980.000 ;
    RECT 497.700 1.400 498.540 980.000 ;
    RECT 498.820 1.400 499.660 980.000 ;
    RECT 499.940 1.400 500.780 980.000 ;
    RECT 501.060 1.400 501.900 980.000 ;
    RECT 502.180 1.400 503.020 980.000 ;
    RECT 503.300 1.400 504.140 980.000 ;
    RECT 504.420 1.400 505.260 980.000 ;
    RECT 505.540 1.400 506.380 980.000 ;
    RECT 506.660 1.400 507.500 980.000 ;
    RECT 507.780 1.400 508.620 980.000 ;
    RECT 508.900 1.400 509.740 980.000 ;
    RECT 510.020 1.400 510.860 980.000 ;
    RECT 511.140 1.400 511.980 980.000 ;
    RECT 512.260 1.400 513.100 980.000 ;
    RECT 513.380 1.400 514.220 980.000 ;
    RECT 514.500 1.400 515.340 980.000 ;
    RECT 515.620 1.400 516.460 980.000 ;
    RECT 516.740 1.400 517.580 980.000 ;
    RECT 517.860 1.400 518.700 980.000 ;
    RECT 518.980 1.400 519.820 980.000 ;
    RECT 520.100 1.400 520.940 980.000 ;
    RECT 521.220 1.400 522.060 980.000 ;
    RECT 522.340 1.400 523.180 980.000 ;
    RECT 523.460 1.400 524.300 980.000 ;
    RECT 524.580 1.400 525.420 980.000 ;
    RECT 525.700 1.400 526.540 980.000 ;
    RECT 526.820 1.400 527.660 980.000 ;
    RECT 527.940 1.400 528.780 980.000 ;
    RECT 529.060 1.400 529.900 980.000 ;
    RECT 530.180 1.400 531.020 980.000 ;
    RECT 531.300 1.400 532.140 980.000 ;
    RECT 532.420 1.400 533.260 980.000 ;
    RECT 533.540 1.400 534.380 980.000 ;
    RECT 534.660 1.400 535.500 980.000 ;
    RECT 535.780 1.400 536.620 980.000 ;
    RECT 536.900 1.400 537.740 980.000 ;
    RECT 538.020 1.400 538.860 980.000 ;
    RECT 539.140 1.400 539.980 980.000 ;
    RECT 540.260 1.400 541.100 980.000 ;
    RECT 541.380 1.400 542.220 980.000 ;
    RECT 542.500 1.400 543.340 980.000 ;
    RECT 543.620 1.400 544.460 980.000 ;
    RECT 544.740 1.400 545.580 980.000 ;
    RECT 545.860 1.400 546.700 980.000 ;
    RECT 546.980 1.400 547.820 980.000 ;
    RECT 548.100 1.400 548.940 980.000 ;
    RECT 549.220 1.400 550.060 980.000 ;
    RECT 550.340 1.400 551.180 980.000 ;
    RECT 551.460 1.400 552.300 980.000 ;
    RECT 552.580 1.400 553.420 980.000 ;
    RECT 553.700 1.400 554.540 980.000 ;
    RECT 554.820 1.400 555.660 980.000 ;
    RECT 555.940 1.400 556.780 980.000 ;
    RECT 557.060 1.400 557.900 980.000 ;
    RECT 558.180 1.400 559.020 980.000 ;
    RECT 559.300 1.400 560.140 980.000 ;
    RECT 560.420 1.400 561.260 980.000 ;
    RECT 561.540 1.400 562.380 980.000 ;
    RECT 562.660 1.400 563.500 980.000 ;
    RECT 563.780 1.400 564.620 980.000 ;
    RECT 564.900 1.400 565.740 980.000 ;
    RECT 566.020 1.400 566.860 980.000 ;
    RECT 567.140 1.400 567.980 980.000 ;
    RECT 568.260 1.400 569.100 980.000 ;
    RECT 569.380 1.400 570.220 980.000 ;
    RECT 570.500 1.400 571.340 980.000 ;
    RECT 571.620 1.400 572.460 980.000 ;
    RECT 572.740 1.400 573.580 980.000 ;
    RECT 573.860 1.400 574.700 980.000 ;
    RECT 574.980 1.400 575.820 980.000 ;
    RECT 576.100 1.400 576.940 980.000 ;
    RECT 577.220 1.400 578.060 980.000 ;
    RECT 578.340 1.400 579.180 980.000 ;
    RECT 579.460 1.400 580.300 980.000 ;
    RECT 580.580 1.400 581.420 980.000 ;
    RECT 581.700 1.400 582.540 980.000 ;
    RECT 582.820 1.400 583.660 980.000 ;
    RECT 583.940 1.400 584.780 980.000 ;
    RECT 585.060 1.400 585.900 980.000 ;
    RECT 586.180 1.400 587.020 980.000 ;
    RECT 587.300 1.400 588.140 980.000 ;
    RECT 588.420 1.400 589.260 980.000 ;
    RECT 589.540 1.400 590.380 980.000 ;
    RECT 590.660 1.400 591.500 980.000 ;
    RECT 591.780 1.400 592.620 980.000 ;
    RECT 592.900 1.400 593.740 980.000 ;
    RECT 594.020 1.400 594.860 980.000 ;
    RECT 595.140 1.400 595.980 980.000 ;
    RECT 596.260 1.400 597.100 980.000 ;
    RECT 597.380 1.400 598.220 980.000 ;
    RECT 598.500 1.400 599.340 980.000 ;
    RECT 599.620 1.400 600.460 980.000 ;
    RECT 600.740 1.400 601.580 980.000 ;
    RECT 601.860 1.400 602.700 980.000 ;
    RECT 602.980 1.400 603.820 980.000 ;
    RECT 604.100 1.400 604.940 980.000 ;
    RECT 605.220 1.400 606.060 980.000 ;
    RECT 606.340 1.400 607.180 980.000 ;
    RECT 607.460 1.400 608.300 980.000 ;
    RECT 608.580 1.400 609.420 980.000 ;
    RECT 609.700 1.400 610.540 980.000 ;
    RECT 610.820 1.400 611.660 980.000 ;
    RECT 611.940 1.400 612.780 980.000 ;
    RECT 613.060 1.400 613.900 980.000 ;
    RECT 614.180 1.400 615.020 980.000 ;
    RECT 615.300 1.400 616.140 980.000 ;
    RECT 616.420 1.400 617.260 980.000 ;
    RECT 617.540 1.400 618.380 980.000 ;
    RECT 618.660 1.400 619.500 980.000 ;
    RECT 619.780 1.400 620.620 980.000 ;
    RECT 620.900 1.400 621.740 980.000 ;
    RECT 622.020 1.400 622.860 980.000 ;
    RECT 623.140 1.400 623.980 980.000 ;
    RECT 624.260 1.400 625.100 980.000 ;
    RECT 625.380 1.400 626.220 980.000 ;
    RECT 626.500 1.400 627.340 980.000 ;
    RECT 627.620 1.400 628.460 980.000 ;
    RECT 628.740 1.400 629.580 980.000 ;
    RECT 629.860 1.400 630.700 980.000 ;
    RECT 630.980 1.400 631.820 980.000 ;
    RECT 632.100 1.400 632.940 980.000 ;
    RECT 633.220 1.400 634.060 980.000 ;
    RECT 634.340 1.400 635.180 980.000 ;
    RECT 635.460 1.400 636.300 980.000 ;
    RECT 636.580 1.400 637.420 980.000 ;
    RECT 637.700 1.400 638.540 980.000 ;
    RECT 638.820 1.400 639.660 980.000 ;
    RECT 639.940 1.400 640.780 980.000 ;
    RECT 641.060 1.400 641.900 980.000 ;
    RECT 642.180 1.400 643.020 980.000 ;
    RECT 643.300 1.400 644.140 980.000 ;
    RECT 644.420 1.400 645.260 980.000 ;
    RECT 645.540 1.400 646.380 980.000 ;
    RECT 646.660 1.400 647.500 980.000 ;
    RECT 647.780 1.400 648.620 980.000 ;
    RECT 648.900 1.400 649.740 980.000 ;
    RECT 650.020 1.400 650.860 980.000 ;
    RECT 651.140 1.400 651.980 980.000 ;
    RECT 652.260 1.400 653.100 980.000 ;
    RECT 653.380 1.400 654.220 980.000 ;
    RECT 654.500 1.400 655.340 980.000 ;
    RECT 655.620 1.400 656.460 980.000 ;
    RECT 656.740 1.400 657.580 980.000 ;
    RECT 657.860 1.400 658.700 980.000 ;
    RECT 658.980 1.400 659.820 980.000 ;
    RECT 660.100 1.400 660.940 980.000 ;
    RECT 661.220 1.400 662.060 980.000 ;
    RECT 662.340 1.400 663.180 980.000 ;
    RECT 663.460 1.400 664.300 980.000 ;
    RECT 664.580 1.400 665.420 980.000 ;
    RECT 665.700 1.400 666.540 980.000 ;
    RECT 666.820 1.400 667.660 980.000 ;
    RECT 667.940 1.400 668.780 980.000 ;
    RECT 669.060 1.400 669.900 980.000 ;
    RECT 670.180 1.400 671.020 980.000 ;
    RECT 671.300 1.400 672.140 980.000 ;
    RECT 672.420 1.400 673.260 980.000 ;
    RECT 673.540 1.400 674.380 980.000 ;
    RECT 674.660 1.400 675.500 980.000 ;
    RECT 675.780 1.400 676.620 980.000 ;
    RECT 676.900 1.400 677.740 980.000 ;
    RECT 678.020 1.400 678.860 980.000 ;
    RECT 679.140 1.400 679.980 980.000 ;
    RECT 680.260 1.400 681.100 980.000 ;
    RECT 681.380 1.400 682.220 980.000 ;
    RECT 682.500 1.400 683.340 980.000 ;
    RECT 683.620 1.400 684.460 980.000 ;
    RECT 684.740 1.400 685.580 980.000 ;
    RECT 685.860 1.400 686.700 980.000 ;
    RECT 686.980 1.400 687.820 980.000 ;
    RECT 688.100 1.400 688.940 980.000 ;
    RECT 689.220 1.400 690.060 980.000 ;
    RECT 690.340 1.400 691.180 980.000 ;
    RECT 691.460 1.400 692.300 980.000 ;
    RECT 692.580 1.400 693.420 980.000 ;
    RECT 693.700 1.400 694.540 980.000 ;
    RECT 694.820 1.400 695.660 980.000 ;
    RECT 695.940 1.400 696.780 980.000 ;
    RECT 697.060 1.400 697.900 980.000 ;
    RECT 698.180 1.400 699.020 980.000 ;
    RECT 699.300 1.400 700.140 980.000 ;
    RECT 700.420 1.400 701.260 980.000 ;
    RECT 701.540 1.400 702.380 980.000 ;
    RECT 702.660 1.400 703.500 980.000 ;
    RECT 703.780 1.400 704.620 980.000 ;
    RECT 704.900 1.400 705.740 980.000 ;
    RECT 706.020 1.400 706.860 980.000 ;
    RECT 707.140 1.400 707.980 980.000 ;
    RECT 708.260 1.400 709.100 980.000 ;
    RECT 709.380 1.400 710.220 980.000 ;
    RECT 710.500 1.400 711.340 980.000 ;
    RECT 711.620 1.400 712.460 980.000 ;
    RECT 712.740 1.400 713.580 980.000 ;
    RECT 713.860 1.400 714.700 980.000 ;
    RECT 714.980 1.400 715.820 980.000 ;
    RECT 716.100 1.400 716.940 980.000 ;
    RECT 717.220 1.400 718.060 980.000 ;
    RECT 718.340 1.400 719.180 980.000 ;
    RECT 719.460 1.400 720.300 980.000 ;
    RECT 720.580 1.400 721.420 980.000 ;
    RECT 721.700 1.400 722.540 980.000 ;
    RECT 722.820 1.400 723.660 980.000 ;
    RECT 723.940 1.400 724.780 980.000 ;
    RECT 725.060 1.400 725.900 980.000 ;
    RECT 726.180 1.400 727.020 980.000 ;
    RECT 727.300 1.400 728.140 980.000 ;
    RECT 728.420 1.400 729.260 980.000 ;
    RECT 729.540 1.400 730.380 980.000 ;
    RECT 730.660 1.400 731.500 980.000 ;
    RECT 731.780 1.400 732.620 980.000 ;
    RECT 732.900 1.400 733.740 980.000 ;
    RECT 734.020 1.400 734.860 980.000 ;
    RECT 735.140 1.400 735.980 980.000 ;
    RECT 736.260 1.400 737.100 980.000 ;
    RECT 737.380 1.400 738.220 980.000 ;
    RECT 738.500 1.400 739.340 980.000 ;
    RECT 739.620 1.400 740.460 980.000 ;
    RECT 740.740 1.400 741.580 980.000 ;
    RECT 741.860 1.400 742.700 980.000 ;
    RECT 742.980 1.400 743.820 980.000 ;
    RECT 744.100 1.400 744.940 980.000 ;
    RECT 745.220 1.400 746.060 980.000 ;
    RECT 746.340 1.400 747.180 980.000 ;
    RECT 747.460 1.400 748.300 980.000 ;
    RECT 748.580 1.400 749.420 980.000 ;
    RECT 749.700 1.400 750.540 980.000 ;
    RECT 750.820 1.400 751.660 980.000 ;
    RECT 751.940 1.400 752.780 980.000 ;
    RECT 753.060 1.400 753.900 980.000 ;
    RECT 754.180 1.400 755.020 980.000 ;
    RECT 755.300 1.400 756.140 980.000 ;
    RECT 756.420 1.400 757.260 980.000 ;
    RECT 757.540 1.400 758.380 980.000 ;
    RECT 758.660 1.400 759.500 980.000 ;
    RECT 759.780 1.400 760.620 980.000 ;
    RECT 760.900 1.400 761.740 980.000 ;
    RECT 762.020 1.400 762.860 980.000 ;
    RECT 763.140 1.400 763.980 980.000 ;
    RECT 764.260 1.400 765.100 980.000 ;
    RECT 765.380 1.400 766.220 980.000 ;
    RECT 766.500 1.400 767.340 980.000 ;
    RECT 767.620 1.400 768.460 980.000 ;
    RECT 768.740 1.400 769.580 980.000 ;
    RECT 769.860 1.400 770.700 980.000 ;
    RECT 770.980 1.400 771.820 980.000 ;
    RECT 772.100 1.400 772.940 980.000 ;
    RECT 773.220 1.400 774.060 980.000 ;
    RECT 774.340 1.400 775.180 980.000 ;
    RECT 775.460 1.400 776.300 980.000 ;
    RECT 776.580 1.400 777.420 980.000 ;
    RECT 777.700 1.400 778.540 980.000 ;
    RECT 778.820 1.400 779.660 980.000 ;
    RECT 779.940 1.400 780.780 980.000 ;
    RECT 781.060 1.400 781.900 980.000 ;
    RECT 782.180 1.400 783.020 980.000 ;
    RECT 783.300 1.400 784.140 980.000 ;
    RECT 784.420 1.400 785.260 980.000 ;
    RECT 785.540 1.400 786.380 980.000 ;
    RECT 786.660 1.400 787.500 980.000 ;
    RECT 787.780 1.400 788.620 980.000 ;
    RECT 788.900 1.400 789.740 980.000 ;
    RECT 790.020 1.400 790.860 980.000 ;
    RECT 791.140 1.400 791.980 980.000 ;
    RECT 792.260 1.400 793.100 980.000 ;
    RECT 793.380 1.400 794.220 980.000 ;
    RECT 794.500 1.400 795.340 980.000 ;
    RECT 795.620 1.400 796.460 980.000 ;
    RECT 796.740 1.400 797.580 980.000 ;
    RECT 797.860 1.400 798.700 980.000 ;
    RECT 798.980 1.400 799.820 980.000 ;
    RECT 800.100 1.400 800.940 980.000 ;
    RECT 801.220 1.400 802.060 980.000 ;
    RECT 802.340 1.400 803.180 980.000 ;
    RECT 803.460 1.400 804.300 980.000 ;
    RECT 804.580 1.400 805.420 980.000 ;
    RECT 805.700 1.400 806.540 980.000 ;
    RECT 806.820 1.400 807.660 980.000 ;
    RECT 807.940 1.400 808.780 980.000 ;
    RECT 809.060 1.400 809.900 980.000 ;
    RECT 810.180 1.400 811.020 980.000 ;
    RECT 811.300 1.400 812.140 980.000 ;
    RECT 812.420 1.400 813.260 980.000 ;
    RECT 813.540 1.400 814.380 980.000 ;
    RECT 814.660 1.400 815.500 980.000 ;
    RECT 815.780 1.400 816.620 980.000 ;
    RECT 816.900 1.400 817.740 980.000 ;
    RECT 818.020 1.400 818.860 980.000 ;
    RECT 819.140 1.400 819.980 980.000 ;
    RECT 820.260 1.400 821.100 980.000 ;
    RECT 821.380 1.400 822.220 980.000 ;
    RECT 822.500 1.400 823.340 980.000 ;
    RECT 823.620 1.400 824.460 980.000 ;
    RECT 824.740 1.400 825.580 980.000 ;
    RECT 825.860 1.400 826.700 980.000 ;
    RECT 826.980 1.400 827.820 980.000 ;
    RECT 828.100 1.400 828.940 980.000 ;
    RECT 829.220 1.400 830.060 980.000 ;
    RECT 830.340 1.400 831.180 980.000 ;
    RECT 831.460 1.400 832.300 980.000 ;
    RECT 832.580 1.400 833.420 980.000 ;
    RECT 833.700 1.400 834.540 980.000 ;
    RECT 834.820 1.400 835.660 980.000 ;
    RECT 835.940 1.400 836.780 980.000 ;
    RECT 837.060 1.400 837.900 980.000 ;
    RECT 838.180 1.400 839.020 980.000 ;
    RECT 839.300 1.400 840.140 980.000 ;
    RECT 840.420 1.400 841.260 980.000 ;
    RECT 841.540 1.400 842.380 980.000 ;
    RECT 842.660 1.400 843.500 980.000 ;
    RECT 843.780 1.400 844.620 980.000 ;
    RECT 844.900 1.400 845.740 980.000 ;
    RECT 846.020 1.400 846.860 980.000 ;
    RECT 847.140 1.400 847.980 980.000 ;
    RECT 848.260 1.400 849.100 980.000 ;
    RECT 849.380 1.400 850.220 980.000 ;
    RECT 850.500 1.400 851.340 980.000 ;
    RECT 851.620 1.400 852.460 980.000 ;
    RECT 852.740 1.400 853.580 980.000 ;
    RECT 853.860 1.400 854.700 980.000 ;
    RECT 854.980 1.400 855.820 980.000 ;
    RECT 856.100 1.400 856.940 980.000 ;
    RECT 857.220 1.400 858.060 980.000 ;
    RECT 858.340 1.400 859.180 980.000 ;
    RECT 859.460 1.400 860.300 980.000 ;
    RECT 860.580 1.400 861.420 980.000 ;
    RECT 861.700 1.400 862.540 980.000 ;
    RECT 862.820 1.400 863.660 980.000 ;
    RECT 863.940 1.400 864.780 980.000 ;
    RECT 865.060 1.400 865.900 980.000 ;
    RECT 866.180 1.400 867.020 980.000 ;
    RECT 867.300 1.400 868.140 980.000 ;
    RECT 868.420 1.400 869.260 980.000 ;
    RECT 869.540 1.400 870.380 980.000 ;
    RECT 870.660 1.400 871.500 980.000 ;
    RECT 871.780 1.400 872.620 980.000 ;
    RECT 872.900 1.400 873.740 980.000 ;
    RECT 874.020 1.400 874.860 980.000 ;
    RECT 875.140 1.400 875.980 980.000 ;
    RECT 876.260 1.400 877.100 980.000 ;
    RECT 877.380 1.400 878.220 980.000 ;
    RECT 878.500 1.400 879.340 980.000 ;
    RECT 879.620 1.400 880.460 980.000 ;
    RECT 880.740 1.400 881.580 980.000 ;
    RECT 881.860 1.400 882.700 980.000 ;
    RECT 882.980 1.400 883.820 980.000 ;
    RECT 884.100 1.400 884.940 980.000 ;
    RECT 885.220 1.400 886.060 980.000 ;
    RECT 886.340 1.400 887.180 980.000 ;
    RECT 887.460 1.400 888.300 980.000 ;
    RECT 888.580 1.400 889.420 980.000 ;
    RECT 889.700 1.400 890.540 980.000 ;
    RECT 890.820 1.400 891.660 980.000 ;
    RECT 891.940 1.400 892.780 980.000 ;
    RECT 893.060 1.400 893.900 980.000 ;
    RECT 894.180 1.400 895.020 980.000 ;
    RECT 895.300 1.400 896.140 980.000 ;
    RECT 896.420 1.400 897.260 980.000 ;
    RECT 897.540 1.400 898.380 980.000 ;
    RECT 898.660 1.400 899.500 980.000 ;
    RECT 899.780 1.400 900.620 980.000 ;
    RECT 900.900 1.400 901.740 980.000 ;
    RECT 902.020 1.400 902.860 980.000 ;
    RECT 903.140 1.400 903.980 980.000 ;
    RECT 904.260 1.400 905.100 980.000 ;
    RECT 905.380 1.400 906.220 980.000 ;
    RECT 906.500 1.400 907.340 980.000 ;
    RECT 907.620 1.400 908.460 980.000 ;
    RECT 908.740 1.400 909.580 980.000 ;
    RECT 909.860 1.400 910.700 980.000 ;
    RECT 910.980 1.400 911.820 980.000 ;
    RECT 912.100 1.400 912.940 980.000 ;
    RECT 913.220 1.400 914.060 980.000 ;
    RECT 914.340 1.400 915.180 980.000 ;
    RECT 915.460 1.400 916.300 980.000 ;
    RECT 916.580 1.400 917.420 980.000 ;
    RECT 917.700 1.400 918.540 980.000 ;
    RECT 918.820 1.400 919.660 980.000 ;
    RECT 919.940 1.400 920.780 980.000 ;
    RECT 921.060 1.400 921.900 980.000 ;
    RECT 922.180 1.400 923.020 980.000 ;
    RECT 923.300 1.400 924.140 980.000 ;
    RECT 924.420 1.400 925.260 980.000 ;
    RECT 925.540 1.400 926.380 980.000 ;
    RECT 926.660 1.400 927.500 980.000 ;
    RECT 927.780 1.400 928.620 980.000 ;
    RECT 928.900 1.400 929.740 980.000 ;
    RECT 930.020 1.400 930.860 980.000 ;
    RECT 931.140 1.400 931.980 980.000 ;
    RECT 932.260 1.400 933.100 980.000 ;
    RECT 933.380 1.400 934.220 980.000 ;
    RECT 934.500 1.400 935.340 980.000 ;
    RECT 935.620 1.400 936.460 980.000 ;
    RECT 936.740 1.400 937.580 980.000 ;
    RECT 937.860 1.400 938.700 980.000 ;
    RECT 938.980 1.400 939.820 980.000 ;
    RECT 940.100 1.400 940.940 980.000 ;
    RECT 941.220 1.400 942.060 980.000 ;
    RECT 942.340 1.400 943.180 980.000 ;
    RECT 943.460 1.400 944.300 980.000 ;
    RECT 944.580 1.400 945.420 980.000 ;
    RECT 945.700 1.400 946.540 980.000 ;
    RECT 946.820 1.400 947.660 980.000 ;
    RECT 947.940 1.400 948.780 980.000 ;
    RECT 949.060 1.400 949.900 980.000 ;
    RECT 950.180 1.400 951.020 980.000 ;
    RECT 951.300 1.400 952.140 980.000 ;
    RECT 952.420 1.400 953.260 980.000 ;
    RECT 953.540 1.400 954.380 980.000 ;
    RECT 954.660 1.400 955.500 980.000 ;
    RECT 955.780 1.400 956.620 980.000 ;
    RECT 956.900 1.400 957.740 980.000 ;
    RECT 958.020 1.400 958.860 980.000 ;
    RECT 959.140 1.400 959.980 980.000 ;
    RECT 960.260 1.400 961.100 980.000 ;
    RECT 961.380 1.400 962.220 980.000 ;
    RECT 962.500 1.400 963.340 980.000 ;
    RECT 963.620 1.400 964.460 980.000 ;
    RECT 964.740 1.400 965.580 980.000 ;
    RECT 965.860 1.400 966.700 980.000 ;
    RECT 966.980 1.400 967.820 980.000 ;
    RECT 968.100 1.400 968.940 980.000 ;
    RECT 969.220 1.400 970.060 980.000 ;
    RECT 970.340 1.400 971.180 980.000 ;
    RECT 971.460 1.400 972.300 980.000 ;
    RECT 972.580 1.400 973.420 980.000 ;
    RECT 973.700 1.400 974.540 980.000 ;
    RECT 974.820 1.400 975.660 980.000 ;
    RECT 975.940 1.400 976.780 980.000 ;
    RECT 977.060 1.400 977.900 980.000 ;
    RECT 978.180 1.400 979.020 980.000 ;
    RECT 979.300 1.400 980.140 980.000 ;
    RECT 980.420 1.400 981.260 980.000 ;
    RECT 981.540 1.400 982.380 980.000 ;
    RECT 982.660 1.400 983.500 980.000 ;
    RECT 983.780 1.400 984.620 980.000 ;
    RECT 984.900 1.400 985.740 980.000 ;
    RECT 986.020 1.400 986.860 980.000 ;
    RECT 987.140 1.400 987.980 980.000 ;
    RECT 988.260 1.400 989.100 980.000 ;
    RECT 989.380 1.400 990.220 980.000 ;
    RECT 990.500 1.400 991.340 980.000 ;
    RECT 991.620 1.400 992.460 980.000 ;
    RECT 992.740 1.400 993.580 980.000 ;
    RECT 993.860 1.400 994.700 980.000 ;
    RECT 994.980 1.400 995.820 980.000 ;
    RECT 996.100 1.400 996.940 980.000 ;
    RECT 997.220 1.400 998.060 980.000 ;
    RECT 998.340 1.400 999.180 980.000 ;
    RECT 999.460 1.400 1000.300 980.000 ;
    RECT 1000.580 1.400 1001.420 980.000 ;
    RECT 1001.700 1.400 1002.540 980.000 ;
    RECT 1002.820 1.400 1003.660 980.000 ;
    RECT 1003.940 1.400 1004.780 980.000 ;
    RECT 1005.060 1.400 1005.900 980.000 ;
    RECT 1006.180 1.400 1007.020 980.000 ;
    RECT 1007.300 1.400 1008.140 980.000 ;
    RECT 1008.420 1.400 1009.260 980.000 ;
    RECT 1009.540 1.400 1010.380 980.000 ;
    RECT 1010.660 1.400 1011.500 980.000 ;
    RECT 1011.780 1.400 1012.620 980.000 ;
    RECT 1012.900 1.400 1013.740 980.000 ;
    RECT 1014.020 1.400 1014.860 980.000 ;
    RECT 1015.140 1.400 1015.980 980.000 ;
    RECT 1016.260 1.400 1017.100 980.000 ;
    RECT 1017.380 1.400 1018.220 980.000 ;
    RECT 1018.500 1.400 1019.340 980.000 ;
    RECT 1019.620 1.400 1020.460 980.000 ;
    RECT 1020.740 1.400 1021.580 980.000 ;
    RECT 1021.860 1.400 1022.700 980.000 ;
    RECT 1022.980 1.400 1023.820 980.000 ;
    RECT 1024.100 1.400 1024.940 980.000 ;
    RECT 1025.220 1.400 1026.060 980.000 ;
    RECT 1026.340 1.400 1027.180 980.000 ;
    RECT 1027.460 1.400 1028.300 980.000 ;
    RECT 1028.580 1.400 1029.420 980.000 ;
    RECT 1029.700 1.400 1030.540 980.000 ;
    RECT 1030.820 1.400 1031.660 980.000 ;
    RECT 1031.940 1.400 1032.780 980.000 ;
    RECT 1033.060 1.400 1033.900 980.000 ;
    RECT 1034.180 1.400 1035.020 980.000 ;
    RECT 1035.300 1.400 1036.140 980.000 ;
    RECT 1036.420 1.400 1037.260 980.000 ;
    RECT 1037.540 1.400 1038.380 980.000 ;
    RECT 1038.660 1.400 1039.500 980.000 ;
    RECT 1039.780 1.400 1040.620 980.000 ;
    RECT 1040.900 1.400 1041.740 980.000 ;
    RECT 1042.020 1.400 1042.860 980.000 ;
    RECT 1043.140 1.400 1043.980 980.000 ;
    RECT 1044.260 1.400 1045.100 980.000 ;
    RECT 1045.380 1.400 1046.220 980.000 ;
    RECT 1046.500 1.400 1047.340 980.000 ;
    RECT 1047.620 1.400 1048.460 980.000 ;
    RECT 1048.740 1.400 1049.580 980.000 ;
    RECT 1049.860 1.400 1050.700 980.000 ;
    RECT 1050.980 1.400 1051.820 980.000 ;
    RECT 1052.100 1.400 1052.940 980.000 ;
    RECT 1053.220 1.400 1054.060 980.000 ;
    RECT 1054.340 1.400 1055.180 980.000 ;
    RECT 1055.460 1.400 1056.300 980.000 ;
    RECT 1056.580 1.400 1057.420 980.000 ;
    RECT 1057.700 1.400 1058.540 980.000 ;
    RECT 1058.820 1.400 1059.660 980.000 ;
    RECT 1059.940 1.400 1060.780 980.000 ;
    RECT 1061.060 1.400 1061.900 980.000 ;
    RECT 1062.180 1.400 1063.020 980.000 ;
    RECT 1063.300 1.400 1064.140 980.000 ;
    RECT 1064.420 1.400 1065.260 980.000 ;
    RECT 1065.540 1.400 1066.380 980.000 ;
    RECT 1066.660 1.400 1067.500 980.000 ;
    RECT 1067.780 1.400 1068.620 980.000 ;
    RECT 1068.900 1.400 1069.740 980.000 ;
    RECT 1070.020 1.400 1070.860 980.000 ;
    RECT 1071.140 1.400 1071.980 980.000 ;
    RECT 1072.260 1.400 1073.100 980.000 ;
    RECT 1073.380 1.400 1074.220 980.000 ;
    RECT 1074.500 1.400 1075.340 980.000 ;
    RECT 1075.620 1.400 1076.460 980.000 ;
    RECT 1076.740 1.400 1077.580 980.000 ;
    RECT 1077.860 1.400 1078.700 980.000 ;
    RECT 1078.980 1.400 1079.820 980.000 ;
    RECT 1080.100 1.400 1080.940 980.000 ;
    RECT 1081.220 1.400 1082.060 980.000 ;
    RECT 1082.340 1.400 1083.180 980.000 ;
    RECT 1083.460 1.400 1084.300 980.000 ;
    RECT 1084.580 1.400 1085.420 980.000 ;
    RECT 1085.700 1.400 1086.540 980.000 ;
    RECT 1086.820 1.400 1087.660 980.000 ;
    RECT 1087.940 1.400 1088.780 980.000 ;
    RECT 1089.060 1.400 1089.900 980.000 ;
    RECT 1090.180 1.400 1091.020 980.000 ;
    RECT 1091.300 1.400 1092.140 980.000 ;
    RECT 1092.420 1.400 1093.260 980.000 ;
    RECT 1093.540 1.400 1094.380 980.000 ;
    RECT 1094.660 1.400 1095.500 980.000 ;
    RECT 1095.780 1.400 1096.620 980.000 ;
    RECT 1096.900 1.400 1097.740 980.000 ;
    RECT 1098.020 1.400 1098.860 980.000 ;
    RECT 1099.140 1.400 1099.980 980.000 ;
    RECT 1100.260 1.400 1101.100 980.000 ;
    RECT 1101.380 1.400 1102.220 980.000 ;
    RECT 1102.500 1.400 1103.340 980.000 ;
    RECT 1103.620 1.400 1104.460 980.000 ;
    RECT 1104.740 1.400 1105.580 980.000 ;
    RECT 1105.860 1.400 1106.700 980.000 ;
    RECT 1106.980 1.400 1107.820 980.000 ;
    RECT 1108.100 1.400 1108.940 980.000 ;
    RECT 1109.220 1.400 1110.060 980.000 ;
    RECT 1110.340 1.400 1111.180 980.000 ;
    RECT 1111.460 1.400 1112.300 980.000 ;
    RECT 1112.580 1.400 1113.420 980.000 ;
    RECT 1113.700 1.400 1114.540 980.000 ;
    RECT 1114.820 1.400 1115.660 980.000 ;
    RECT 1115.940 1.400 1116.780 980.000 ;
    RECT 1117.060 1.400 1117.900 980.000 ;
    RECT 1118.180 1.400 1119.020 980.000 ;
    RECT 1119.300 1.400 1120.140 980.000 ;
    RECT 1120.420 1.400 1121.260 980.000 ;
    RECT 1121.540 1.400 1122.380 980.000 ;
    RECT 1122.660 1.400 1123.500 980.000 ;
    RECT 1123.780 1.400 1124.620 980.000 ;
    RECT 1124.900 1.400 1125.740 980.000 ;
    RECT 1126.020 1.400 1126.860 980.000 ;
    RECT 1127.140 1.400 1127.980 980.000 ;
    RECT 1128.260 1.400 1129.100 980.000 ;
    RECT 1129.380 1.400 1130.220 980.000 ;
    RECT 1130.500 1.400 1131.340 980.000 ;
    RECT 1131.620 1.400 1132.460 980.000 ;
    RECT 1132.740 1.400 1133.580 980.000 ;
    RECT 1133.860 1.400 1134.700 980.000 ;
    RECT 1134.980 1.400 1135.820 980.000 ;
    RECT 1136.100 1.400 1136.940 980.000 ;
    RECT 1137.220 1.400 1138.060 980.000 ;
    RECT 1138.340 1.400 1139.180 980.000 ;
    RECT 1139.460 1.400 1140.300 980.000 ;
    RECT 1140.580 1.400 1141.420 980.000 ;
    RECT 1141.700 1.400 1142.540 980.000 ;
    RECT 1142.820 1.400 1143.660 980.000 ;
    RECT 1143.940 1.400 1144.780 980.000 ;
    RECT 1145.060 1.400 1145.900 980.000 ;
    RECT 1146.180 1.400 1147.020 980.000 ;
    RECT 1147.300 1.400 1148.140 980.000 ;
    RECT 1148.420 1.400 1149.260 980.000 ;
    RECT 1149.540 1.400 1150.380 980.000 ;
    RECT 1150.660 1.400 1151.500 980.000 ;
    RECT 1151.780 1.400 1152.620 980.000 ;
    RECT 1152.900 1.400 1153.740 980.000 ;
    RECT 1154.020 1.400 1154.860 980.000 ;
    RECT 1155.140 1.400 1155.980 980.000 ;
    RECT 1156.260 1.400 1157.100 980.000 ;
    RECT 1157.380 1.400 1158.220 980.000 ;
    RECT 1158.500 1.400 1159.340 980.000 ;
    RECT 1159.620 1.400 1160.460 980.000 ;
    RECT 1160.740 1.400 1161.580 980.000 ;
    RECT 1161.860 1.400 1162.700 980.000 ;
    RECT 1162.980 1.400 1163.820 980.000 ;
    RECT 1164.100 1.400 1164.940 980.000 ;
    RECT 1165.220 1.400 1166.060 980.000 ;
    RECT 1166.340 1.400 1167.180 980.000 ;
    RECT 1167.460 1.400 1168.300 980.000 ;
    RECT 1168.580 1.400 1169.420 980.000 ;
    RECT 1169.700 1.400 1170.540 980.000 ;
    RECT 1170.820 1.400 1171.660 980.000 ;
    RECT 1171.940 1.400 1172.780 980.000 ;
    RECT 1173.060 1.400 1173.900 980.000 ;
    RECT 1174.180 1.400 1175.020 980.000 ;
    RECT 1175.300 1.400 1176.140 980.000 ;
    RECT 1176.420 1.400 1177.260 980.000 ;
    RECT 1177.540 1.400 1178.380 980.000 ;
    RECT 1178.660 1.400 1179.500 980.000 ;
    RECT 1179.780 1.400 1180.620 980.000 ;
    RECT 1180.900 1.400 1181.740 980.000 ;
    RECT 1182.020 1.400 1182.860 980.000 ;
    RECT 1183.140 1.400 1183.980 980.000 ;
    RECT 1184.260 1.400 1185.100 980.000 ;
    RECT 1185.380 1.400 1186.220 980.000 ;
    RECT 1186.500 1.400 1187.340 980.000 ;
    RECT 1187.620 1.400 1188.460 980.000 ;
    RECT 1188.740 1.400 1189.580 980.000 ;
    RECT 1189.860 1.400 1190.700 980.000 ;
    RECT 1190.980 1.400 1191.820 980.000 ;
    RECT 1192.100 1.400 1192.940 980.000 ;
    RECT 1193.220 1.400 1194.060 980.000 ;
    RECT 1194.340 1.400 1195.180 980.000 ;
    RECT 1195.460 1.400 1196.300 980.000 ;
    RECT 1196.580 1.400 1197.420 980.000 ;
    RECT 1197.700 1.400 1198.540 980.000 ;
    RECT 1198.820 1.400 1199.660 980.000 ;
    RECT 1199.940 1.400 1200.780 980.000 ;
    RECT 1201.060 1.400 1201.900 980.000 ;
    RECT 1202.180 1.400 1203.020 980.000 ;
    RECT 1203.300 1.400 1204.140 980.000 ;
    RECT 1204.420 1.400 1205.260 980.000 ;
    RECT 1205.540 1.400 1206.380 980.000 ;
    RECT 1206.660 1.400 1207.500 980.000 ;
    RECT 1207.780 1.400 1208.620 980.000 ;
    RECT 1208.900 1.400 1209.740 980.000 ;
    RECT 1210.020 1.400 1210.860 980.000 ;
    RECT 1211.140 1.400 1211.980 980.000 ;
    RECT 1212.260 1.400 1213.100 980.000 ;
    RECT 1213.380 1.400 1214.220 980.000 ;
    RECT 1214.500 1.400 1215.340 980.000 ;
    RECT 1215.620 1.400 1216.460 980.000 ;
    RECT 1216.740 1.400 1217.580 980.000 ;
    RECT 1217.860 1.400 1218.700 980.000 ;
    RECT 1218.980 1.400 1219.820 980.000 ;
    RECT 1220.100 1.400 1220.940 980.000 ;
    RECT 1221.220 1.400 1222.060 980.000 ;
    RECT 1222.340 1.400 1223.180 980.000 ;
    RECT 1223.460 1.400 1224.300 980.000 ;
    RECT 1224.580 1.400 1225.420 980.000 ;
    RECT 1225.700 1.400 1226.540 980.000 ;
    RECT 1226.820 1.400 1227.660 980.000 ;
    RECT 1227.940 1.400 1228.780 980.000 ;
    RECT 1229.060 1.400 1229.900 980.000 ;
    RECT 1230.180 1.400 1231.020 980.000 ;
    RECT 1231.300 1.400 1232.140 980.000 ;
    RECT 1232.420 1.400 1233.260 980.000 ;
    RECT 1233.540 1.400 1234.380 980.000 ;
    RECT 1234.660 1.400 1235.500 980.000 ;
    RECT 1235.780 1.400 1236.620 980.000 ;
    RECT 1236.900 1.400 1237.740 980.000 ;
    RECT 1238.020 1.400 1238.860 980.000 ;
    RECT 1239.140 1.400 1239.980 980.000 ;
    RECT 1240.260 1.400 1241.100 980.000 ;
    RECT 1241.380 1.400 1242.220 980.000 ;
    RECT 1242.500 1.400 1243.340 980.000 ;
    RECT 1243.620 1.400 1244.460 980.000 ;
    RECT 1244.740 1.400 1245.580 980.000 ;
    RECT 1245.860 1.400 1246.700 980.000 ;
    RECT 1246.980 1.400 1247.820 980.000 ;
    RECT 1248.100 1.400 1248.940 980.000 ;
    RECT 1249.220 1.400 1250.060 980.000 ;
    RECT 1250.340 1.400 1251.180 980.000 ;
    RECT 1251.460 1.400 1252.300 980.000 ;
    RECT 1252.580 1.400 1253.420 980.000 ;
    RECT 1253.700 1.400 1254.540 980.000 ;
    RECT 1254.820 1.400 1255.660 980.000 ;
    RECT 1255.940 1.400 1256.780 980.000 ;
    RECT 1257.060 1.400 1257.900 980.000 ;
    RECT 1258.180 1.400 1259.020 980.000 ;
    RECT 1259.300 1.400 1260.140 980.000 ;
    RECT 1260.420 1.400 1261.260 980.000 ;
    RECT 1261.540 1.400 1262.380 980.000 ;
    RECT 1262.660 1.400 1263.500 980.000 ;
    RECT 1263.780 1.400 1264.620 980.000 ;
    RECT 1264.900 1.400 1265.740 980.000 ;
    RECT 1266.020 1.400 1266.860 980.000 ;
    RECT 1267.140 1.400 1267.980 980.000 ;
    RECT 1268.260 1.400 1269.100 980.000 ;
    RECT 1269.380 1.400 1270.220 980.000 ;
    RECT 1270.500 1.400 1271.340 980.000 ;
    RECT 1271.620 1.400 1272.460 980.000 ;
    RECT 1272.740 1.400 1273.580 980.000 ;
    RECT 1273.860 1.400 1274.700 980.000 ;
    RECT 1274.980 1.400 1275.820 980.000 ;
    RECT 1276.100 1.400 1276.940 980.000 ;
    RECT 1277.220 1.400 1278.060 980.000 ;
    RECT 1278.340 1.400 1279.180 980.000 ;
    RECT 1279.460 1.400 1280.300 980.000 ;
    RECT 1280.580 1.400 1281.420 980.000 ;
    RECT 1281.700 1.400 1282.540 980.000 ;
    RECT 1282.820 1.400 1283.660 980.000 ;
    RECT 1283.940 1.400 1284.780 980.000 ;
    RECT 1285.060 1.400 1285.900 980.000 ;
    RECT 1286.180 1.400 1287.020 980.000 ;
    RECT 1287.300 1.400 1288.140 980.000 ;
    RECT 1288.420 1.400 1289.260 980.000 ;
    RECT 1289.540 1.400 1290.380 980.000 ;
    RECT 1290.660 1.400 1291.500 980.000 ;
    RECT 1291.780 1.400 1292.620 980.000 ;
    RECT 1292.900 1.400 1293.740 980.000 ;
    RECT 1294.020 1.400 1294.860 980.000 ;
    RECT 1295.140 1.400 1295.980 980.000 ;
    RECT 1296.260 1.400 1297.100 980.000 ;
    RECT 1297.380 1.400 1298.220 980.000 ;
    RECT 1298.500 1.400 1299.340 980.000 ;
    RECT 1299.620 1.400 1300.460 980.000 ;
    RECT 1300.740 1.400 1301.580 980.000 ;
    RECT 1301.860 1.400 1302.700 980.000 ;
    RECT 1302.980 1.400 1303.820 980.000 ;
    RECT 1304.100 1.400 1304.940 980.000 ;
    RECT 1305.220 1.400 1306.060 980.000 ;
    RECT 1306.340 1.400 1307.180 980.000 ;
    RECT 1307.460 1.400 1308.300 980.000 ;
    RECT 1308.580 1.400 1309.420 980.000 ;
    RECT 1309.700 1.400 1310.540 980.000 ;
    RECT 1310.820 1.400 1311.660 980.000 ;
    RECT 1311.940 1.400 1312.780 980.000 ;
    RECT 1313.060 1.400 1313.900 980.000 ;
    RECT 1314.180 1.400 1315.020 980.000 ;
    RECT 1315.300 1.400 1316.140 980.000 ;
    RECT 1316.420 1.400 1317.260 980.000 ;
    RECT 1317.540 1.400 1318.380 980.000 ;
    RECT 1318.660 1.400 1319.500 980.000 ;
    RECT 1319.780 1.400 1320.620 980.000 ;
    RECT 1320.900 1.400 1321.740 980.000 ;
    RECT 1322.020 1.400 1322.860 980.000 ;
    RECT 1323.140 1.400 1323.980 980.000 ;
    RECT 1324.260 1.400 1325.100 980.000 ;
    RECT 1325.380 1.400 1326.220 980.000 ;
    RECT 1326.500 1.400 1327.340 980.000 ;
    RECT 1327.620 1.400 1328.460 980.000 ;
    RECT 1328.740 1.400 1329.580 980.000 ;
    RECT 1329.860 1.400 1330.700 980.000 ;
    RECT 1330.980 1.400 1331.820 980.000 ;
    RECT 1332.100 1.400 1332.940 980.000 ;
    RECT 1333.220 1.400 1334.060 980.000 ;
    RECT 1334.340 1.400 1335.180 980.000 ;
    RECT 1335.460 1.400 1336.300 980.000 ;
    RECT 1336.580 1.400 1337.420 980.000 ;
    RECT 1337.700 1.400 1338.540 980.000 ;
    RECT 1338.820 1.400 1339.660 980.000 ;
    RECT 1339.940 1.400 1340.780 980.000 ;
    RECT 1341.060 1.400 1341.900 980.000 ;
    RECT 1342.180 1.400 1343.020 980.000 ;
    RECT 1343.300 1.400 1344.140 980.000 ;
    RECT 1344.420 1.400 1345.260 980.000 ;
    RECT 1345.540 1.400 1346.380 980.000 ;
    RECT 1346.660 1.400 1347.500 980.000 ;
    RECT 1347.780 1.400 1348.620 980.000 ;
    RECT 1348.900 1.400 1349.740 980.000 ;
    RECT 1350.020 1.400 1350.860 980.000 ;
    RECT 1351.140 1.400 1351.980 980.000 ;
    RECT 1352.260 1.400 1353.100 980.000 ;
    RECT 1353.380 1.400 1354.220 980.000 ;
    RECT 1354.500 1.400 1355.340 980.000 ;
    RECT 1355.620 1.400 1356.460 980.000 ;
    RECT 1356.740 1.400 1357.580 980.000 ;
    RECT 1357.860 1.400 1358.700 980.000 ;
    RECT 1358.980 1.400 1359.820 980.000 ;
    RECT 1360.100 1.400 1360.940 980.000 ;
    RECT 1361.220 1.400 1362.060 980.000 ;
    RECT 1362.340 1.400 1363.180 980.000 ;
    RECT 1363.460 1.400 1364.300 980.000 ;
    RECT 1364.580 1.400 1365.420 980.000 ;
    RECT 1365.700 1.400 1366.540 980.000 ;
    RECT 1366.820 1.400 1367.660 980.000 ;
    RECT 1367.940 1.400 1368.780 980.000 ;
    RECT 1369.060 1.400 1369.900 980.000 ;
    RECT 1370.180 1.400 1371.020 980.000 ;
    RECT 1371.300 1.400 1372.140 980.000 ;
    RECT 1372.420 1.400 1373.260 980.000 ;
    RECT 1373.540 1.400 1374.380 980.000 ;
    RECT 1374.660 1.400 1375.500 980.000 ;
    RECT 1375.780 1.400 1376.620 980.000 ;
    RECT 1376.900 1.400 1377.740 980.000 ;
    RECT 1378.020 1.400 1378.860 980.000 ;
    RECT 1379.140 1.400 1379.980 980.000 ;
    RECT 1380.260 1.400 1381.100 980.000 ;
    RECT 1381.380 1.400 1382.220 980.000 ;
    RECT 1382.500 1.400 1383.340 980.000 ;
    RECT 1383.620 1.400 1384.460 980.000 ;
    RECT 1384.740 1.400 1385.580 980.000 ;
    RECT 1385.860 1.400 1386.700 980.000 ;
    RECT 1386.980 1.400 1387.820 980.000 ;
    RECT 1388.100 1.400 1388.940 980.000 ;
    RECT 1389.220 1.400 1390.060 980.000 ;
    RECT 1390.340 1.400 1391.180 980.000 ;
    RECT 1391.460 1.400 1392.300 980.000 ;
    RECT 1392.580 1.400 1393.420 980.000 ;
    RECT 1393.700 1.400 1394.540 980.000 ;
    RECT 1394.820 1.400 1395.660 980.000 ;
    RECT 1395.940 1.400 1396.780 980.000 ;
    RECT 1397.060 1.400 1397.900 980.000 ;
    RECT 1398.180 1.400 1399.020 980.000 ;
    RECT 1399.300 1.400 1400.140 980.000 ;
    RECT 1400.420 1.400 1401.260 980.000 ;
    RECT 1401.540 1.400 1402.380 980.000 ;
    RECT 1402.660 1.400 1403.500 980.000 ;
    RECT 1403.780 1.400 1404.620 980.000 ;
    RECT 1404.900 1.400 1405.740 980.000 ;
    RECT 1406.020 1.400 1406.860 980.000 ;
    RECT 1407.140 1.400 1407.980 980.000 ;
    RECT 1408.260 1.400 1409.100 980.000 ;
    RECT 1409.380 1.400 1410.220 980.000 ;
    RECT 1410.500 1.400 1411.340 980.000 ;
    RECT 1411.620 1.400 1412.460 980.000 ;
    RECT 1412.740 1.400 1413.580 980.000 ;
    RECT 1413.860 1.400 1414.700 980.000 ;
    RECT 1414.980 1.400 1415.820 980.000 ;
    RECT 1416.100 1.400 1416.940 980.000 ;
    RECT 1417.220 1.400 1418.060 980.000 ;
    RECT 1418.340 1.400 1419.180 980.000 ;
    RECT 1419.460 1.400 1420.300 980.000 ;
    RECT 1420.580 1.400 1421.420 980.000 ;
    RECT 1421.700 1.400 1422.540 980.000 ;
    RECT 1422.820 1.400 1423.660 980.000 ;
    RECT 1423.940 1.400 1424.780 980.000 ;
    RECT 1425.060 1.400 1425.900 980.000 ;
    RECT 1426.180 1.400 1427.020 980.000 ;
    RECT 1427.300 1.400 1428.140 980.000 ;
    RECT 1428.420 1.400 1429.260 980.000 ;
    RECT 1429.540 1.400 1430.380 980.000 ;
    RECT 1430.660 1.400 1431.500 980.000 ;
    RECT 1431.780 1.400 1432.620 980.000 ;
    RECT 1432.900 1.400 1433.740 980.000 ;
    RECT 1434.020 1.400 1434.860 980.000 ;
    RECT 1435.140 1.400 1435.980 980.000 ;
    RECT 1436.260 1.400 1437.100 980.000 ;
    RECT 1437.380 1.400 1438.220 980.000 ;
    RECT 1438.500 1.400 1439.340 980.000 ;
    RECT 1439.620 1.400 1440.460 980.000 ;
    RECT 1440.740 1.400 1441.580 980.000 ;
    RECT 1441.860 1.400 1442.700 980.000 ;
    RECT 1442.980 1.400 1443.820 980.000 ;
    RECT 1444.100 1.400 1444.940 980.000 ;
    RECT 1445.220 1.400 1446.060 980.000 ;
    RECT 1446.340 1.400 1447.180 980.000 ;
    RECT 1447.460 1.400 1448.300 980.000 ;
    RECT 1448.580 1.400 1449.420 980.000 ;
    RECT 1449.700 1.400 1450.540 980.000 ;
    RECT 1450.820 1.400 1451.660 980.000 ;
    RECT 1451.940 1.400 1452.780 980.000 ;
    RECT 1453.060 1.400 1453.900 980.000 ;
    RECT 1454.180 1.400 1455.020 980.000 ;
    RECT 1455.300 1.400 1456.140 980.000 ;
    RECT 1456.420 1.400 1457.260 980.000 ;
    RECT 1457.540 1.400 1458.380 980.000 ;
    RECT 1458.660 1.400 1459.500 980.000 ;
    RECT 1459.780 1.400 1460.620 980.000 ;
    RECT 1460.900 1.400 1461.740 980.000 ;
    RECT 1462.020 1.400 1462.860 980.000 ;
    RECT 1463.140 1.400 1463.980 980.000 ;
    RECT 1464.260 1.400 1465.100 980.000 ;
    RECT 1465.380 1.400 1466.220 980.000 ;
    RECT 1466.500 1.400 1467.340 980.000 ;
    RECT 1467.620 1.400 1468.460 980.000 ;
    RECT 1468.740 1.400 1469.580 980.000 ;
    RECT 1469.860 1.400 1470.700 980.000 ;
    RECT 1470.980 1.400 1471.820 980.000 ;
    RECT 1472.100 1.400 1472.940 980.000 ;
    RECT 1473.220 1.400 1474.060 980.000 ;
    RECT 1474.340 1.400 1475.180 980.000 ;
    RECT 1475.460 1.400 1476.300 980.000 ;
    RECT 1476.580 1.400 1477.420 980.000 ;
    RECT 1477.700 1.400 1478.540 980.000 ;
    RECT 1478.820 1.400 1479.660 980.000 ;
    RECT 1479.940 1.400 1480.780 980.000 ;
    RECT 1481.060 1.400 1481.900 980.000 ;
    RECT 1482.180 1.400 1483.020 980.000 ;
    RECT 1483.300 1.400 1484.140 980.000 ;
    RECT 1484.420 1.400 1485.260 980.000 ;
    RECT 1485.540 1.400 1486.380 980.000 ;
    RECT 1486.660 1.400 1487.500 980.000 ;
    RECT 1487.780 1.400 1488.620 980.000 ;
    RECT 1488.900 1.400 1489.740 980.000 ;
    RECT 1490.020 1.400 1490.860 980.000 ;
    RECT 1491.140 1.400 1491.980 980.000 ;
    RECT 1492.260 1.400 1493.100 980.000 ;
    RECT 1493.380 1.400 1494.220 980.000 ;
    RECT 1494.500 1.400 1495.340 980.000 ;
    RECT 1495.620 1.400 1496.460 980.000 ;
    RECT 1496.740 1.400 1497.580 980.000 ;
    RECT 1497.860 1.400 1498.700 980.000 ;
    RECT 1498.980 1.400 1499.820 980.000 ;
    RECT 1500.100 1.400 1500.940 980.000 ;
    RECT 1501.220 1.400 1502.060 980.000 ;
    RECT 1502.340 1.400 1503.180 980.000 ;
    RECT 1503.460 1.400 1504.300 980.000 ;
    RECT 1504.580 1.400 1505.420 980.000 ;
    RECT 1505.700 1.400 1506.540 980.000 ;
    RECT 1506.820 1.400 1507.660 980.000 ;
    RECT 1507.940 1.400 1508.780 980.000 ;
    RECT 1509.060 1.400 1509.900 980.000 ;
    RECT 1510.180 1.400 1511.020 980.000 ;
    RECT 1511.300 1.400 1512.140 980.000 ;
    RECT 1512.420 1.400 1513.260 980.000 ;
    RECT 1513.540 1.400 1514.380 980.000 ;
    RECT 1514.660 1.400 1515.500 980.000 ;
    RECT 1515.780 1.400 1516.620 980.000 ;
    RECT 1516.900 1.400 1517.740 980.000 ;
    RECT 1518.020 1.400 1518.860 980.000 ;
    RECT 1519.140 1.400 1519.980 980.000 ;
    RECT 1520.260 1.400 1521.100 980.000 ;
    RECT 1521.380 1.400 1522.220 980.000 ;
    RECT 1522.500 1.400 1523.340 980.000 ;
    RECT 1523.620 1.400 1524.460 980.000 ;
    RECT 1524.740 1.400 1525.580 980.000 ;
    RECT 1525.860 1.400 1526.700 980.000 ;
    RECT 1526.980 1.400 1527.820 980.000 ;
    RECT 1528.100 1.400 1528.940 980.000 ;
    RECT 1529.220 1.400 1530.060 980.000 ;
    RECT 1530.340 1.400 1531.180 980.000 ;
    RECT 1531.460 1.400 1532.300 980.000 ;
    RECT 1532.580 1.400 1533.420 980.000 ;
    RECT 1533.700 1.400 1534.540 980.000 ;
    RECT 1534.820 1.400 1535.660 980.000 ;
    RECT 1535.940 1.400 1536.780 980.000 ;
    RECT 1537.060 1.400 1537.900 980.000 ;
    RECT 1538.180 1.400 1539.020 980.000 ;
    RECT 1539.300 1.400 1540.140 980.000 ;
    RECT 1540.420 1.400 1541.260 980.000 ;
    RECT 1541.540 1.400 1542.380 980.000 ;
    RECT 1542.660 1.400 1543.500 980.000 ;
    RECT 1543.780 1.400 1544.620 980.000 ;
    RECT 1544.900 1.400 1545.740 980.000 ;
    RECT 1546.020 1.400 1546.860 980.000 ;
    RECT 1547.140 1.400 1547.980 980.000 ;
    RECT 1548.260 1.400 1549.100 980.000 ;
    RECT 1549.380 1.400 1550.220 980.000 ;
    RECT 1550.500 1.400 1551.340 980.000 ;
    RECT 1551.620 1.400 1552.460 980.000 ;
    RECT 1552.740 1.400 1553.580 980.000 ;
    RECT 1553.860 1.400 1554.700 980.000 ;
    RECT 1554.980 1.400 1555.820 980.000 ;
    RECT 1556.100 1.400 1556.940 980.000 ;
    RECT 1557.220 1.400 1558.060 980.000 ;
    RECT 1558.340 1.400 1559.180 980.000 ;
    RECT 1559.460 1.400 1560.300 980.000 ;
    RECT 1560.580 1.400 1561.420 980.000 ;
    RECT 1561.700 1.400 1562.540 980.000 ;
    RECT 1562.820 1.400 1563.660 980.000 ;
    RECT 1563.940 1.400 1564.780 980.000 ;
    RECT 1565.060 1.400 1565.900 980.000 ;
    RECT 1566.180 1.400 1567.020 980.000 ;
    RECT 1567.300 1.400 1568.140 980.000 ;
    RECT 1568.420 1.400 1569.260 980.000 ;
    RECT 1569.540 1.400 1570.380 980.000 ;
    RECT 1570.660 1.400 1571.500 980.000 ;
    RECT 1571.780 1.400 1572.620 980.000 ;
    RECT 1572.900 1.400 1573.740 980.000 ;
    RECT 1574.020 1.400 1574.860 980.000 ;
    RECT 1575.140 1.400 1575.980 980.000 ;
    RECT 1576.260 1.400 1577.100 980.000 ;
    RECT 1577.380 1.400 1578.220 980.000 ;
    RECT 1578.500 1.400 1579.340 980.000 ;
    RECT 1579.620 1.400 1580.460 980.000 ;
    RECT 1580.740 1.400 1581.580 980.000 ;
    RECT 1581.860 1.400 1582.700 980.000 ;
    RECT 1582.980 1.400 1583.820 980.000 ;
    RECT 1584.100 1.400 1584.940 980.000 ;
    RECT 1585.220 1.400 1586.060 980.000 ;
    RECT 1586.340 1.400 1587.180 980.000 ;
    RECT 1587.460 1.400 1588.300 980.000 ;
    RECT 1588.580 1.400 1589.420 980.000 ;
    RECT 1589.700 1.400 1590.540 980.000 ;
    RECT 1590.820 1.400 1591.660 980.000 ;
    RECT 1591.940 1.400 1592.780 980.000 ;
    RECT 1593.060 1.400 1593.900 980.000 ;
    RECT 1594.180 1.400 1595.020 980.000 ;
    RECT 1595.300 1.400 1596.140 980.000 ;
    RECT 1596.420 1.400 1597.260 980.000 ;
    RECT 1597.540 1.400 1598.380 980.000 ;
    RECT 1598.660 1.400 1599.500 980.000 ;
    RECT 1599.780 1.400 1600.620 980.000 ;
    RECT 1600.900 1.400 1601.740 980.000 ;
    RECT 1602.020 1.400 1602.860 980.000 ;
    RECT 1603.140 1.400 1603.980 980.000 ;
    RECT 1604.260 1.400 1605.100 980.000 ;
    RECT 1605.380 1.400 1606.220 980.000 ;
    RECT 1606.500 1.400 1607.340 980.000 ;
    RECT 1607.620 1.400 1608.460 980.000 ;
    RECT 1608.740 1.400 1609.580 980.000 ;
    RECT 1609.860 1.400 1610.700 980.000 ;
    RECT 1610.980 1.400 1611.820 980.000 ;
    RECT 1612.100 1.400 1612.940 980.000 ;
    RECT 1613.220 1.400 1614.060 980.000 ;
    RECT 1614.340 1.400 1615.180 980.000 ;
    RECT 1615.460 1.400 1616.300 980.000 ;
    RECT 1616.580 1.400 1617.420 980.000 ;
    RECT 1617.700 1.400 1618.540 980.000 ;
    RECT 1618.820 1.400 1619.660 980.000 ;
    RECT 1619.940 1.400 1620.780 980.000 ;
    RECT 1621.060 1.400 1621.900 980.000 ;
    RECT 1622.180 1.400 1623.020 980.000 ;
    RECT 1623.300 1.400 1624.140 980.000 ;
    RECT 1624.420 1.400 1625.260 980.000 ;
    RECT 1625.540 1.400 1626.380 980.000 ;
    RECT 1626.660 1.400 1627.500 980.000 ;
    RECT 1627.780 1.400 1628.620 980.000 ;
    RECT 1628.900 1.400 1629.740 980.000 ;
    RECT 1630.020 1.400 1630.860 980.000 ;
    RECT 1631.140 1.400 1631.980 980.000 ;
    RECT 1632.260 1.400 1633.100 980.000 ;
    RECT 1633.380 1.400 1634.220 980.000 ;
    RECT 1634.500 1.400 1635.340 980.000 ;
    RECT 1635.620 1.400 1636.460 980.000 ;
    RECT 1636.740 1.400 1637.580 980.000 ;
    RECT 1637.860 1.400 1638.700 980.000 ;
    RECT 1638.980 1.400 1639.820 980.000 ;
    RECT 1640.100 1.400 1640.940 980.000 ;
    RECT 1641.220 1.400 1642.060 980.000 ;
    RECT 1642.340 1.400 1643.180 980.000 ;
    RECT 1643.460 1.400 1644.300 980.000 ;
    RECT 1644.580 1.400 1645.420 980.000 ;
    RECT 1645.700 1.400 1646.540 980.000 ;
    RECT 1646.820 1.400 1647.660 980.000 ;
    RECT 1647.940 1.400 1648.780 980.000 ;
    RECT 1649.060 1.400 1649.900 980.000 ;
    RECT 1650.180 1.400 1651.020 980.000 ;
    RECT 1651.300 1.400 1652.140 980.000 ;
    RECT 1652.420 1.400 1653.260 980.000 ;
    RECT 1653.540 1.400 1654.380 980.000 ;
    RECT 1654.660 1.400 1655.500 980.000 ;
    RECT 1655.780 1.400 1656.620 980.000 ;
    RECT 1656.900 1.400 1657.740 980.000 ;
    RECT 1658.020 1.400 1658.860 980.000 ;
    RECT 1659.140 1.400 1659.980 980.000 ;
    RECT 1660.260 1.400 1661.100 980.000 ;
    RECT 1661.380 1.400 1662.220 980.000 ;
    RECT 1662.500 1.400 1663.340 980.000 ;
    RECT 1663.620 1.400 1664.460 980.000 ;
    RECT 1664.740 1.400 1665.580 980.000 ;
    RECT 1665.860 1.400 1666.700 980.000 ;
    RECT 1666.980 1.400 1667.820 980.000 ;
    RECT 1668.100 1.400 1668.940 980.000 ;
    RECT 1669.220 1.400 1670.060 980.000 ;
    RECT 1670.340 1.400 1671.180 980.000 ;
    RECT 1671.460 1.400 1672.300 980.000 ;
    RECT 1672.580 1.400 1673.420 980.000 ;
    RECT 1673.700 1.400 1674.540 980.000 ;
    RECT 1674.820 1.400 1675.660 980.000 ;
    RECT 1675.940 1.400 1676.780 980.000 ;
    RECT 1677.060 1.400 1677.900 980.000 ;
    RECT 1678.180 1.400 1679.020 980.000 ;
    RECT 1679.300 1.400 1680.140 980.000 ;
    RECT 1680.420 1.400 1681.260 980.000 ;
    RECT 1681.540 1.400 1682.380 980.000 ;
    RECT 1682.660 1.400 1683.500 980.000 ;
    RECT 1683.780 1.400 1684.620 980.000 ;
    RECT 1684.900 1.400 1685.740 980.000 ;
    RECT 1686.020 1.400 1686.860 980.000 ;
    RECT 1687.140 1.400 1687.980 980.000 ;
    RECT 1688.260 1.400 1689.100 980.000 ;
    RECT 1689.380 1.400 1690.220 980.000 ;
    RECT 1690.500 1.400 1691.340 980.000 ;
    RECT 1691.620 1.400 1692.460 980.000 ;
    RECT 1692.740 1.400 1693.580 980.000 ;
    RECT 1693.860 1.400 1694.700 980.000 ;
    RECT 1694.980 1.400 1695.820 980.000 ;
    RECT 1696.100 1.400 1696.940 980.000 ;
    RECT 1697.220 1.400 1698.060 980.000 ;
    RECT 1698.340 1.400 1699.180 980.000 ;
    RECT 1699.460 1.400 1700.300 980.000 ;
    RECT 1700.580 1.400 1701.420 980.000 ;
    RECT 1701.700 1.400 1702.540 980.000 ;
    RECT 1702.820 1.400 1703.660 980.000 ;
    RECT 1703.940 1.400 1704.780 980.000 ;
    RECT 1705.060 1.400 1705.900 980.000 ;
    RECT 1706.180 1.400 1707.020 980.000 ;
    RECT 1707.300 1.400 1708.140 980.000 ;
    RECT 1708.420 1.400 1709.260 980.000 ;
    RECT 1709.540 1.400 1710.380 980.000 ;
    RECT 1710.660 1.400 1711.500 980.000 ;
    RECT 1711.780 1.400 1712.620 980.000 ;
    RECT 1712.900 1.400 1713.740 980.000 ;
    RECT 1714.020 1.400 1714.860 980.000 ;
    RECT 1715.140 1.400 1715.980 980.000 ;
    RECT 1716.260 1.400 1717.100 980.000 ;
    RECT 1717.380 1.400 1718.220 980.000 ;
    RECT 1718.500 1.400 1719.340 980.000 ;
    RECT 1719.620 1.400 1720.460 980.000 ;
    RECT 1720.740 1.400 1721.580 980.000 ;
    RECT 1721.860 1.400 1722.700 980.000 ;
    RECT 1722.980 1.400 1723.820 980.000 ;
    RECT 1724.100 1.400 1724.940 980.000 ;
    RECT 1725.220 1.400 1726.060 980.000 ;
    RECT 1726.340 1.400 1727.180 980.000 ;
    RECT 1727.460 1.400 1728.300 980.000 ;
    RECT 1728.580 1.400 1729.420 980.000 ;
    RECT 1729.700 1.400 1730.540 980.000 ;
    RECT 1730.820 1.400 1731.660 980.000 ;
    RECT 1731.940 1.400 1732.780 980.000 ;
    RECT 1733.060 1.400 1733.900 980.000 ;
    RECT 1734.180 1.400 1735.020 980.000 ;
    RECT 1735.300 1.400 1736.140 980.000 ;
    RECT 1736.420 1.400 1737.260 980.000 ;
    RECT 1737.540 1.400 1738.380 980.000 ;
    RECT 1738.660 1.400 1739.500 980.000 ;
    RECT 1739.780 1.400 1740.620 980.000 ;
    RECT 1740.900 1.400 1741.740 980.000 ;
    RECT 1742.020 1.400 1742.860 980.000 ;
    RECT 1743.140 1.400 1743.980 980.000 ;
    RECT 1744.260 1.400 1745.100 980.000 ;
    RECT 1745.380 1.400 1746.220 980.000 ;
    RECT 1746.500 1.400 1747.340 980.000 ;
    RECT 1747.620 1.400 1748.460 980.000 ;
    RECT 1748.740 1.400 1749.580 980.000 ;
    RECT 1749.860 1.400 1750.700 980.000 ;
    RECT 1750.980 1.400 1751.820 980.000 ;
    RECT 1752.100 1.400 1752.940 980.000 ;
    RECT 1753.220 1.400 1754.060 980.000 ;
    RECT 1754.340 1.400 1755.180 980.000 ;
    RECT 1755.460 1.400 1756.300 980.000 ;
    RECT 1756.580 1.400 1757.420 980.000 ;
    RECT 1757.700 1.400 1758.540 980.000 ;
    RECT 1758.820 1.400 1759.660 980.000 ;
    RECT 1759.940 1.400 1760.780 980.000 ;
    RECT 1761.060 1.400 1761.900 980.000 ;
    RECT 1762.180 1.400 1763.020 980.000 ;
    RECT 1763.300 1.400 1764.140 980.000 ;
    RECT 1764.420 1.400 1765.260 980.000 ;
    RECT 1765.540 1.400 1766.380 980.000 ;
    RECT 1766.660 1.400 1767.500 980.000 ;
    RECT 1767.780 1.400 1768.620 980.000 ;
    RECT 1768.900 1.400 1769.740 980.000 ;
    RECT 1770.020 1.400 1770.860 980.000 ;
    RECT 1771.140 1.400 1771.980 980.000 ;
    RECT 1772.260 1.400 1773.100 980.000 ;
    RECT 1773.380 1.400 1774.220 980.000 ;
    RECT 1774.500 1.400 1775.340 980.000 ;
    RECT 1775.620 1.400 1776.460 980.000 ;
    RECT 1776.740 1.400 1777.580 980.000 ;
    RECT 1777.860 1.400 1778.700 980.000 ;
    RECT 1778.980 1.400 1779.820 980.000 ;
    RECT 1780.100 1.400 1780.940 980.000 ;
    RECT 1781.220 1.400 1782.060 980.000 ;
    RECT 1782.340 1.400 1783.180 980.000 ;
    RECT 1783.460 1.400 1784.300 980.000 ;
    RECT 1784.580 1.400 1785.420 980.000 ;
    RECT 1785.700 1.400 1786.540 980.000 ;
    RECT 1786.820 1.400 1787.660 980.000 ;
    RECT 1787.940 1.400 1788.780 980.000 ;
    RECT 1789.060 1.400 1789.900 980.000 ;
    RECT 1790.180 1.400 1791.020 980.000 ;
    RECT 1791.300 1.400 1792.140 980.000 ;
    RECT 1792.420 1.400 1793.260 980.000 ;
    RECT 1793.540 1.400 1794.380 980.000 ;
    RECT 1794.660 1.400 1795.500 980.000 ;
    RECT 1795.780 1.400 1796.620 980.000 ;
    RECT 1796.900 1.400 1797.740 980.000 ;
    RECT 1798.020 1.400 1798.860 980.000 ;
    RECT 1799.140 1.400 1799.980 980.000 ;
    RECT 1800.260 1.400 1801.100 980.000 ;
    RECT 1801.380 1.400 1802.220 980.000 ;
    RECT 1802.500 1.400 1803.340 980.000 ;
    RECT 1803.620 1.400 1804.460 980.000 ;
    RECT 1804.740 1.400 1805.580 980.000 ;
    RECT 1805.860 1.400 1806.700 980.000 ;
    RECT 1806.980 1.400 1807.820 980.000 ;
    RECT 1808.100 1.400 1808.940 980.000 ;
    RECT 1809.220 1.400 1810.060 980.000 ;
    RECT 1810.340 1.400 1811.180 980.000 ;
    RECT 1811.460 1.400 1812.300 980.000 ;
    RECT 1812.580 1.400 1813.420 980.000 ;
    RECT 1813.700 1.400 1814.540 980.000 ;
    RECT 1814.820 1.400 1815.660 980.000 ;
    RECT 1815.940 1.400 1816.780 980.000 ;
    RECT 1817.060 1.400 1817.900 980.000 ;
    RECT 1818.180 1.400 1819.020 980.000 ;
    RECT 1819.300 1.400 1820.140 980.000 ;
    RECT 1820.420 1.400 1821.260 980.000 ;
    RECT 1821.540 1.400 1822.380 980.000 ;
    RECT 1822.660 1.400 1823.500 980.000 ;
    RECT 1823.780 1.400 1824.620 980.000 ;
    RECT 1824.900 1.400 1825.740 980.000 ;
    RECT 1826.020 1.400 1826.860 980.000 ;
    RECT 1827.140 1.400 1827.980 980.000 ;
    RECT 1828.260 1.400 1829.100 980.000 ;
    RECT 1829.380 1.400 1830.220 980.000 ;
    RECT 1830.500 1.400 1832.740 980.000 ;
    LAYER OVERLAP ;
    RECT 0 0 1832.740 981.400 ;
  END
END sram_512x1024_1r1w

END LIBRARY
