VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_32x128_2r1w
  FOREIGN fakeram_32x128_2r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 96.710 BY 250.600 ;
  CLASS BLOCK ;
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 0.805 0.140 0.875 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.140 13.895 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.140 26.915 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.140 39.935 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.140 52.955 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.905 0.140 65.975 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.140 78.995 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.945 0.140 92.015 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 0.805 96.710 0.875 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 13.825 96.710 13.895 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 26.845 96.710 26.915 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 39.865 96.710 39.935 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 52.885 96.710 52.955 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 65.905 96.710 65.975 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 78.925 96.710 78.995 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 91.945 96.710 92.015 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1.105 0.000 1.175 0.140 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 3.005 0.000 3.075 0.140 ;
    END
  END w0_wd_in[17]
  PIN w0_wd_in[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 4.905 0.000 4.975 0.140 ;
    END
  END w0_wd_in[18]
  PIN w0_wd_in[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 6.805 0.000 6.875 0.140 ;
    END
  END w0_wd_in[19]
  PIN w0_wd_in[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 8.705 0.000 8.775 0.140 ;
    END
  END w0_wd_in[20]
  PIN w0_wd_in[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 10.605 0.000 10.675 0.140 ;
    END
  END w0_wd_in[21]
  PIN w0_wd_in[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 12.505 0.000 12.575 0.140 ;
    END
  END w0_wd_in[22]
  PIN w0_wd_in[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 14.405 0.000 14.475 0.140 ;
    END
  END w0_wd_in[23]
  PIN w0_wd_in[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 16.305 0.000 16.375 0.140 ;
    END
  END w0_wd_in[24]
  PIN w0_wd_in[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 18.205 0.000 18.275 0.140 ;
    END
  END w0_wd_in[25]
  PIN w0_wd_in[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 20.105 0.000 20.175 0.140 ;
    END
  END w0_wd_in[26]
  PIN w0_wd_in[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 22.005 0.000 22.075 0.140 ;
    END
  END w0_wd_in[27]
  PIN w0_wd_in[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 23.905 0.000 23.975 0.140 ;
    END
  END w0_wd_in[28]
  PIN w0_wd_in[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 25.805 0.000 25.875 0.140 ;
    END
  END w0_wd_in[29]
  PIN w0_wd_in[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 27.705 0.000 27.775 0.140 ;
    END
  END w0_wd_in[30]
  PIN w0_wd_in[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 29.605 0.000 29.675 0.140 ;
    END
  END w0_wd_in[31]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 31.505 0.000 31.575 0.140 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 33.405 0.000 33.475 0.140 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 35.305 0.000 35.375 0.140 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 37.205 0.000 37.275 0.140 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 39.105 0.000 39.175 0.140 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 41.005 0.000 41.075 0.140 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 42.905 0.000 42.975 0.140 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 44.805 0.000 44.875 0.140 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 46.705 0.000 46.775 0.140 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 48.605 0.000 48.675 0.140 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 50.505 0.000 50.575 0.140 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 52.405 0.000 52.475 0.140 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 54.305 0.000 54.375 0.140 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 56.205 0.000 56.275 0.140 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 58.105 0.000 58.175 0.140 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 60.005 0.000 60.075 0.140 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1.105 250.460 1.175 250.600 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 3.385 250.460 3.455 250.600 ;
    END
  END r0_rd_out[17]
  PIN r0_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 5.665 250.460 5.735 250.600 ;
    END
  END r0_rd_out[18]
  PIN r0_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 7.945 250.460 8.015 250.600 ;
    END
  END r0_rd_out[19]
  PIN r0_rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 10.225 250.460 10.295 250.600 ;
    END
  END r0_rd_out[20]
  PIN r0_rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 12.505 250.460 12.575 250.600 ;
    END
  END r0_rd_out[21]
  PIN r0_rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 14.785 250.460 14.855 250.600 ;
    END
  END r0_rd_out[22]
  PIN r0_rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 17.065 250.460 17.135 250.600 ;
    END
  END r0_rd_out[23]
  PIN r0_rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 19.345 250.460 19.415 250.600 ;
    END
  END r0_rd_out[24]
  PIN r0_rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 21.625 250.460 21.695 250.600 ;
    END
  END r0_rd_out[25]
  PIN r0_rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 23.905 250.460 23.975 250.600 ;
    END
  END r0_rd_out[26]
  PIN r0_rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 26.185 250.460 26.255 250.600 ;
    END
  END r0_rd_out[27]
  PIN r0_rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 28.465 250.460 28.535 250.600 ;
    END
  END r0_rd_out[28]
  PIN r0_rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 30.745 250.460 30.815 250.600 ;
    END
  END r0_rd_out[29]
  PIN r0_rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 33.025 250.460 33.095 250.600 ;
    END
  END r0_rd_out[30]
  PIN r0_rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 35.305 250.460 35.375 250.600 ;
    END
  END r0_rd_out[31]
  PIN r1_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 61.905 0.000 61.975 0.140 ;
    END
  END r1_rd_out[0]
  PIN r1_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 63.805 0.000 63.875 0.140 ;
    END
  END r1_rd_out[1]
  PIN r1_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 65.705 0.000 65.775 0.140 ;
    END
  END r1_rd_out[2]
  PIN r1_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 67.605 0.000 67.675 0.140 ;
    END
  END r1_rd_out[3]
  PIN r1_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 69.505 0.000 69.575 0.140 ;
    END
  END r1_rd_out[4]
  PIN r1_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 71.405 0.000 71.475 0.140 ;
    END
  END r1_rd_out[5]
  PIN r1_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 73.305 0.000 73.375 0.140 ;
    END
  END r1_rd_out[6]
  PIN r1_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 75.205 0.000 75.275 0.140 ;
    END
  END r1_rd_out[7]
  PIN r1_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 77.105 0.000 77.175 0.140 ;
    END
  END r1_rd_out[8]
  PIN r1_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 79.005 0.000 79.075 0.140 ;
    END
  END r1_rd_out[9]
  PIN r1_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 80.905 0.000 80.975 0.140 ;
    END
  END r1_rd_out[10]
  PIN r1_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 82.805 0.000 82.875 0.140 ;
    END
  END r1_rd_out[11]
  PIN r1_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 84.705 0.000 84.775 0.140 ;
    END
  END r1_rd_out[12]
  PIN r1_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 86.605 0.000 86.675 0.140 ;
    END
  END r1_rd_out[13]
  PIN r1_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 88.505 0.000 88.575 0.140 ;
    END
  END r1_rd_out[14]
  PIN r1_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 90.405 0.000 90.475 0.140 ;
    END
  END r1_rd_out[15]
  PIN r1_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 37.585 250.460 37.655 250.600 ;
    END
  END r1_rd_out[16]
  PIN r1_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 39.865 250.460 39.935 250.600 ;
    END
  END r1_rd_out[17]
  PIN r1_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 42.145 250.460 42.215 250.600 ;
    END
  END r1_rd_out[18]
  PIN r1_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 44.425 250.460 44.495 250.600 ;
    END
  END r1_rd_out[19]
  PIN r1_rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 46.705 250.460 46.775 250.600 ;
    END
  END r1_rd_out[20]
  PIN r1_rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 48.985 250.460 49.055 250.600 ;
    END
  END r1_rd_out[21]
  PIN r1_rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 51.265 250.460 51.335 250.600 ;
    END
  END r1_rd_out[22]
  PIN r1_rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 53.545 250.460 53.615 250.600 ;
    END
  END r1_rd_out[23]
  PIN r1_rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 55.825 250.460 55.895 250.600 ;
    END
  END r1_rd_out[24]
  PIN r1_rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 58.105 250.460 58.175 250.600 ;
    END
  END r1_rd_out[25]
  PIN r1_rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 60.385 250.460 60.455 250.600 ;
    END
  END r1_rd_out[26]
  PIN r1_rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 62.665 250.460 62.735 250.600 ;
    END
  END r1_rd_out[27]
  PIN r1_rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 64.945 250.460 65.015 250.600 ;
    END
  END r1_rd_out[28]
  PIN r1_rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 67.225 250.460 67.295 250.600 ;
    END
  END r1_rd_out[29]
  PIN r1_rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 69.505 250.460 69.575 250.600 ;
    END
  END r1_rd_out[30]
  PIN r1_rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 71.785 250.460 71.855 250.600 ;
    END
  END r1_rd_out[31]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.965 0.140 105.035 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.985 0.140 118.055 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.005 0.140 131.075 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.025 0.140 144.095 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 104.965 96.710 105.035 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 117.985 96.710 118.055 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 131.005 96.710 131.075 ;
    END
  END w0_addr_in[6]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.045 0.140 157.115 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.065 0.140 170.135 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.085 0.140 183.155 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.105 0.140 196.175 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 144.025 96.710 144.095 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 157.045 96.710 157.115 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 170.065 96.710 170.135 ;
    END
  END r0_addr_in[6]
  PIN r1_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.125 0.140 209.195 ;
    END
  END r1_addr_in[0]
  PIN r1_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.145 0.140 222.215 ;
    END
  END r1_addr_in[1]
  PIN r1_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.165 0.140 235.235 ;
    END
  END r1_addr_in[2]
  PIN r1_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.185 0.140 248.255 ;
    END
  END r1_addr_in[3]
  PIN r1_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 183.085 96.710 183.155 ;
    END
  END r1_addr_in[4]
  PIN r1_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 196.105 96.710 196.175 ;
    END
  END r1_addr_in[5]
  PIN r1_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 96.570 209.125 96.710 209.195 ;
    END
  END r1_addr_in[6]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 74.065 250.460 74.135 250.600 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 76.345 250.460 76.415 250.600 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 78.625 250.460 78.695 250.600 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 80.905 250.460 80.975 250.600 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 83.185 250.460 83.255 250.600 ;
    END
  END r0_clk
  PIN r1_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 85.465 250.460 85.535 250.600 ;
    END
  END r1_ce_in
  PIN r1_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 87.745 250.460 87.815 250.600 ;
    END
  END r1_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 0.430 0.700 0.710 249.900 ;
      RECT 2.670 0.700 2.950 249.900 ;
      RECT 4.910 0.700 5.190 249.900 ;
      RECT 7.150 0.700 7.430 249.900 ;
      RECT 9.390 0.700 9.670 249.900 ;
      RECT 11.630 0.700 11.910 249.900 ;
      RECT 13.870 0.700 14.150 249.900 ;
      RECT 16.110 0.700 16.390 249.900 ;
      RECT 18.350 0.700 18.630 249.900 ;
      RECT 20.590 0.700 20.870 249.900 ;
      RECT 22.830 0.700 23.110 249.900 ;
      RECT 25.070 0.700 25.350 249.900 ;
      RECT 27.310 0.700 27.590 249.900 ;
      RECT 29.550 0.700 29.830 249.900 ;
      RECT 31.790 0.700 32.070 249.900 ;
      RECT 34.030 0.700 34.310 249.900 ;
      RECT 36.270 0.700 36.550 249.900 ;
      RECT 38.510 0.700 38.790 249.900 ;
      RECT 40.750 0.700 41.030 249.900 ;
      RECT 42.990 0.700 43.270 249.900 ;
      RECT 45.230 0.700 45.510 249.900 ;
      RECT 47.470 0.700 47.750 249.900 ;
      RECT 49.710 0.700 49.990 249.900 ;
      RECT 51.950 0.700 52.230 249.900 ;
      RECT 54.190 0.700 54.470 249.900 ;
      RECT 56.430 0.700 56.710 249.900 ;
      RECT 58.670 0.700 58.950 249.900 ;
      RECT 60.910 0.700 61.190 249.900 ;
      RECT 63.150 0.700 63.430 249.900 ;
      RECT 65.390 0.700 65.670 249.900 ;
      RECT 67.630 0.700 67.910 249.900 ;
      RECT 69.870 0.700 70.150 249.900 ;
      RECT 72.110 0.700 72.390 249.900 ;
      RECT 74.350 0.700 74.630 249.900 ;
      RECT 76.590 0.700 76.870 249.900 ;
      RECT 78.830 0.700 79.110 249.900 ;
      RECT 81.070 0.700 81.350 249.900 ;
      RECT 83.310 0.700 83.590 249.900 ;
      RECT 85.550 0.700 85.830 249.900 ;
      RECT 87.790 0.700 88.070 249.900 ;
      RECT 90.030 0.700 90.310 249.900 ;
      RECT 92.270 0.700 92.550 249.900 ;
      RECT 94.510 0.700 94.790 249.900 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 0.430 0.700 0.710 249.900 ;
      RECT 2.670 0.700 2.950 249.900 ;
      RECT 4.910 0.700 5.190 249.900 ;
      RECT 7.150 0.700 7.430 249.900 ;
      RECT 9.390 0.700 9.670 249.900 ;
      RECT 11.630 0.700 11.910 249.900 ;
      RECT 13.870 0.700 14.150 249.900 ;
      RECT 16.110 0.700 16.390 249.900 ;
      RECT 18.350 0.700 18.630 249.900 ;
      RECT 20.590 0.700 20.870 249.900 ;
      RECT 22.830 0.700 23.110 249.900 ;
      RECT 25.070 0.700 25.350 249.900 ;
      RECT 27.310 0.700 27.590 249.900 ;
      RECT 29.550 0.700 29.830 249.900 ;
      RECT 31.790 0.700 32.070 249.900 ;
      RECT 34.030 0.700 34.310 249.900 ;
      RECT 36.270 0.700 36.550 249.900 ;
      RECT 38.510 0.700 38.790 249.900 ;
      RECT 40.750 0.700 41.030 249.900 ;
      RECT 42.990 0.700 43.270 249.900 ;
      RECT 45.230 0.700 45.510 249.900 ;
      RECT 47.470 0.700 47.750 249.900 ;
      RECT 49.710 0.700 49.990 249.900 ;
      RECT 51.950 0.700 52.230 249.900 ;
      RECT 54.190 0.700 54.470 249.900 ;
      RECT 56.430 0.700 56.710 249.900 ;
      RECT 58.670 0.700 58.950 249.900 ;
      RECT 60.910 0.700 61.190 249.900 ;
      RECT 63.150 0.700 63.430 249.900 ;
      RECT 65.390 0.700 65.670 249.900 ;
      RECT 67.630 0.700 67.910 249.900 ;
      RECT 69.870 0.700 70.150 249.900 ;
      RECT 72.110 0.700 72.390 249.900 ;
      RECT 74.350 0.700 74.630 249.900 ;
      RECT 76.590 0.700 76.870 249.900 ;
      RECT 78.830 0.700 79.110 249.900 ;
      RECT 81.070 0.700 81.350 249.900 ;
      RECT 83.310 0.700 83.590 249.900 ;
      RECT 85.550 0.700 85.830 249.900 ;
      RECT 87.790 0.700 88.070 249.900 ;
      RECT 90.030 0.700 90.310 249.900 ;
      RECT 92.270 0.700 92.550 249.900 ;
      RECT 94.510 0.700 94.790 249.900 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 96.710 250.600 ;
    LAYER metal2 ;
    RECT 0 0 96.710 250.600 ;
    LAYER metal3 ;
    RECT 0 0 96.710 250.600 ;
    LAYER metal4 ;
    RECT 0 0 96.710 250.600 ;
    LAYER OVERLAP ;
    RECT 0 0 96.710 250.600 ;
  END
END fakeram_32x128_2r1w

END LIBRARY
