VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO liteeth_1rw1r_32w384d_32_sram
  FOREIGN liteeth_1rw1r_32w384d_32_sram 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 568.100 BY 544.000 ;
  CLASS BLOCK ;
  PIN w_mask_rw1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 5.850 0.800 6.150 ;
    END
  END w_mask_rw1[0]
  PIN w_mask_rw1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 10.050 0.800 10.350 ;
    END
  END w_mask_rw1[1]
  PIN w_mask_rw1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.250 0.800 14.550 ;
    END
  END w_mask_rw1[2]
  PIN w_mask_rw1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 18.450 0.800 18.750 ;
    END
  END w_mask_rw1[3]
  PIN w_mask_rw1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.650 0.800 22.950 ;
    END
  END w_mask_rw1[4]
  PIN w_mask_rw1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 26.850 0.800 27.150 ;
    END
  END w_mask_rw1[5]
  PIN w_mask_rw1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.050 0.800 31.350 ;
    END
  END w_mask_rw1[6]
  PIN w_mask_rw1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 35.250 0.800 35.550 ;
    END
  END w_mask_rw1[7]
  PIN w_mask_rw1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.450 0.800 39.750 ;
    END
  END w_mask_rw1[8]
  PIN w_mask_rw1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 43.650 0.800 43.950 ;
    END
  END w_mask_rw1[9]
  PIN w_mask_rw1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 47.850 0.800 48.150 ;
    END
  END w_mask_rw1[10]
  PIN w_mask_rw1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 52.050 0.800 52.350 ;
    END
  END w_mask_rw1[11]
  PIN w_mask_rw1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 56.250 0.800 56.550 ;
    END
  END w_mask_rw1[12]
  PIN w_mask_rw1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 60.450 0.800 60.750 ;
    END
  END w_mask_rw1[13]
  PIN w_mask_rw1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 64.650 0.800 64.950 ;
    END
  END w_mask_rw1[14]
  PIN w_mask_rw1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 68.850 0.800 69.150 ;
    END
  END w_mask_rw1[15]
  PIN w_mask_rw1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 73.050 0.800 73.350 ;
    END
  END w_mask_rw1[16]
  PIN w_mask_rw1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 77.250 0.800 77.550 ;
    END
  END w_mask_rw1[17]
  PIN w_mask_rw1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 81.450 0.800 81.750 ;
    END
  END w_mask_rw1[18]
  PIN w_mask_rw1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 85.650 0.800 85.950 ;
    END
  END w_mask_rw1[19]
  PIN w_mask_rw1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.850 0.800 90.150 ;
    END
  END w_mask_rw1[20]
  PIN w_mask_rw1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 94.050 0.800 94.350 ;
    END
  END w_mask_rw1[21]
  PIN w_mask_rw1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 98.250 0.800 98.550 ;
    END
  END w_mask_rw1[22]
  PIN w_mask_rw1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 102.450 0.800 102.750 ;
    END
  END w_mask_rw1[23]
  PIN w_mask_rw1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 106.650 0.800 106.950 ;
    END
  END w_mask_rw1[24]
  PIN w_mask_rw1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 110.850 0.800 111.150 ;
    END
  END w_mask_rw1[25]
  PIN w_mask_rw1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 115.050 0.800 115.350 ;
    END
  END w_mask_rw1[26]
  PIN w_mask_rw1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 119.250 0.800 119.550 ;
    END
  END w_mask_rw1[27]
  PIN w_mask_rw1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 123.450 0.800 123.750 ;
    END
  END w_mask_rw1[28]
  PIN w_mask_rw1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 127.650 0.800 127.950 ;
    END
  END w_mask_rw1[29]
  PIN w_mask_rw1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 131.850 0.800 132.150 ;
    END
  END w_mask_rw1[30]
  PIN w_mask_rw1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 136.050 0.800 136.350 ;
    END
  END w_mask_rw1[31]
  PIN rd_out_rw1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 140.250 0.800 140.550 ;
    END
  END rd_out_rw1[0]
  PIN rd_out_rw1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 144.450 0.800 144.750 ;
    END
  END rd_out_rw1[1]
  PIN rd_out_rw1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 148.650 0.800 148.950 ;
    END
  END rd_out_rw1[2]
  PIN rd_out_rw1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 152.850 0.800 153.150 ;
    END
  END rd_out_rw1[3]
  PIN rd_out_rw1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 157.050 0.800 157.350 ;
    END
  END rd_out_rw1[4]
  PIN rd_out_rw1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 161.250 0.800 161.550 ;
    END
  END rd_out_rw1[5]
  PIN rd_out_rw1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 165.450 0.800 165.750 ;
    END
  END rd_out_rw1[6]
  PIN rd_out_rw1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 169.650 0.800 169.950 ;
    END
  END rd_out_rw1[7]
  PIN rd_out_rw1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 173.850 0.800 174.150 ;
    END
  END rd_out_rw1[8]
  PIN rd_out_rw1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 178.050 0.800 178.350 ;
    END
  END rd_out_rw1[9]
  PIN rd_out_rw1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 182.250 0.800 182.550 ;
    END
  END rd_out_rw1[10]
  PIN rd_out_rw1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 186.450 0.800 186.750 ;
    END
  END rd_out_rw1[11]
  PIN rd_out_rw1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 190.650 0.800 190.950 ;
    END
  END rd_out_rw1[12]
  PIN rd_out_rw1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 194.850 0.800 195.150 ;
    END
  END rd_out_rw1[13]
  PIN rd_out_rw1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 199.050 0.800 199.350 ;
    END
  END rd_out_rw1[14]
  PIN rd_out_rw1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 203.250 0.800 203.550 ;
    END
  END rd_out_rw1[15]
  PIN rd_out_rw1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 207.450 0.800 207.750 ;
    END
  END rd_out_rw1[16]
  PIN rd_out_rw1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 211.650 0.800 211.950 ;
    END
  END rd_out_rw1[17]
  PIN rd_out_rw1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 215.850 0.800 216.150 ;
    END
  END rd_out_rw1[18]
  PIN rd_out_rw1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 220.050 0.800 220.350 ;
    END
  END rd_out_rw1[19]
  PIN rd_out_rw1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 224.250 0.800 224.550 ;
    END
  END rd_out_rw1[20]
  PIN rd_out_rw1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 228.450 0.800 228.750 ;
    END
  END rd_out_rw1[21]
  PIN rd_out_rw1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 232.650 0.800 232.950 ;
    END
  END rd_out_rw1[22]
  PIN rd_out_rw1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 236.850 0.800 237.150 ;
    END
  END rd_out_rw1[23]
  PIN rd_out_rw1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 241.050 0.800 241.350 ;
    END
  END rd_out_rw1[24]
  PIN rd_out_rw1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 245.250 0.800 245.550 ;
    END
  END rd_out_rw1[25]
  PIN rd_out_rw1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 249.450 0.800 249.750 ;
    END
  END rd_out_rw1[26]
  PIN rd_out_rw1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 253.650 0.800 253.950 ;
    END
  END rd_out_rw1[27]
  PIN rd_out_rw1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 257.850 0.800 258.150 ;
    END
  END rd_out_rw1[28]
  PIN rd_out_rw1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 262.050 0.800 262.350 ;
    END
  END rd_out_rw1[29]
  PIN rd_out_rw1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 266.250 0.800 266.550 ;
    END
  END rd_out_rw1[30]
  PIN rd_out_rw1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 270.450 0.800 270.750 ;
    END
  END rd_out_rw1[31]
  PIN rd_out_r1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 274.650 0.800 274.950 ;
    END
  END rd_out_r1[0]
  PIN rd_out_r1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 278.850 0.800 279.150 ;
    END
  END rd_out_r1[1]
  PIN rd_out_r1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 283.050 0.800 283.350 ;
    END
  END rd_out_r1[2]
  PIN rd_out_r1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 287.250 0.800 287.550 ;
    END
  END rd_out_r1[3]
  PIN rd_out_r1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 291.450 0.800 291.750 ;
    END
  END rd_out_r1[4]
  PIN rd_out_r1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 295.650 0.800 295.950 ;
    END
  END rd_out_r1[5]
  PIN rd_out_r1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 299.850 0.800 300.150 ;
    END
  END rd_out_r1[6]
  PIN rd_out_r1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 304.050 0.800 304.350 ;
    END
  END rd_out_r1[7]
  PIN rd_out_r1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 308.250 0.800 308.550 ;
    END
  END rd_out_r1[8]
  PIN rd_out_r1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 312.450 0.800 312.750 ;
    END
  END rd_out_r1[9]
  PIN rd_out_r1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 316.650 0.800 316.950 ;
    END
  END rd_out_r1[10]
  PIN rd_out_r1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 320.850 0.800 321.150 ;
    END
  END rd_out_r1[11]
  PIN rd_out_r1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 325.050 0.800 325.350 ;
    END
  END rd_out_r1[12]
  PIN rd_out_r1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 329.250 0.800 329.550 ;
    END
  END rd_out_r1[13]
  PIN rd_out_r1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 333.450 0.800 333.750 ;
    END
  END rd_out_r1[14]
  PIN rd_out_r1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 337.650 0.800 337.950 ;
    END
  END rd_out_r1[15]
  PIN rd_out_r1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 341.850 0.800 342.150 ;
    END
  END rd_out_r1[16]
  PIN rd_out_r1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 346.050 0.800 346.350 ;
    END
  END rd_out_r1[17]
  PIN rd_out_r1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 350.250 0.800 350.550 ;
    END
  END rd_out_r1[18]
  PIN rd_out_r1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 354.450 0.800 354.750 ;
    END
  END rd_out_r1[19]
  PIN rd_out_r1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 358.650 0.800 358.950 ;
    END
  END rd_out_r1[20]
  PIN rd_out_r1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 362.850 0.800 363.150 ;
    END
  END rd_out_r1[21]
  PIN rd_out_r1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 367.050 0.800 367.350 ;
    END
  END rd_out_r1[22]
  PIN rd_out_r1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 371.250 0.800 371.550 ;
    END
  END rd_out_r1[23]
  PIN rd_out_r1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 375.450 0.800 375.750 ;
    END
  END rd_out_r1[24]
  PIN rd_out_r1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 379.650 0.800 379.950 ;
    END
  END rd_out_r1[25]
  PIN rd_out_r1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 383.850 0.800 384.150 ;
    END
  END rd_out_r1[26]
  PIN rd_out_r1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 388.050 0.800 388.350 ;
    END
  END rd_out_r1[27]
  PIN rd_out_r1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 392.250 0.800 392.550 ;
    END
  END rd_out_r1[28]
  PIN rd_out_r1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 396.450 0.800 396.750 ;
    END
  END rd_out_r1[29]
  PIN rd_out_r1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 400.650 0.800 400.950 ;
    END
  END rd_out_r1[30]
  PIN rd_out_r1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 404.850 0.800 405.150 ;
    END
  END rd_out_r1[31]
  PIN wd_in_rw1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 409.050 0.800 409.350 ;
    END
  END wd_in_rw1[0]
  PIN wd_in_rw1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 413.250 0.800 413.550 ;
    END
  END wd_in_rw1[1]
  PIN wd_in_rw1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 417.450 0.800 417.750 ;
    END
  END wd_in_rw1[2]
  PIN wd_in_rw1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 421.650 0.800 421.950 ;
    END
  END wd_in_rw1[3]
  PIN wd_in_rw1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 425.850 0.800 426.150 ;
    END
  END wd_in_rw1[4]
  PIN wd_in_rw1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 430.050 0.800 430.350 ;
    END
  END wd_in_rw1[5]
  PIN wd_in_rw1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 434.250 0.800 434.550 ;
    END
  END wd_in_rw1[6]
  PIN wd_in_rw1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 438.450 0.800 438.750 ;
    END
  END wd_in_rw1[7]
  PIN wd_in_rw1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 442.650 0.800 442.950 ;
    END
  END wd_in_rw1[8]
  PIN wd_in_rw1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 446.850 0.800 447.150 ;
    END
  END wd_in_rw1[9]
  PIN wd_in_rw1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 451.050 0.800 451.350 ;
    END
  END wd_in_rw1[10]
  PIN wd_in_rw1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 455.250 0.800 455.550 ;
    END
  END wd_in_rw1[11]
  PIN wd_in_rw1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 459.450 0.800 459.750 ;
    END
  END wd_in_rw1[12]
  PIN wd_in_rw1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 463.650 0.800 463.950 ;
    END
  END wd_in_rw1[13]
  PIN wd_in_rw1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 467.850 0.800 468.150 ;
    END
  END wd_in_rw1[14]
  PIN wd_in_rw1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 472.050 0.800 472.350 ;
    END
  END wd_in_rw1[15]
  PIN wd_in_rw1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 476.250 0.800 476.550 ;
    END
  END wd_in_rw1[16]
  PIN wd_in_rw1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 480.450 0.800 480.750 ;
    END
  END wd_in_rw1[17]
  PIN wd_in_rw1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 484.650 0.800 484.950 ;
    END
  END wd_in_rw1[18]
  PIN wd_in_rw1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 488.850 0.800 489.150 ;
    END
  END wd_in_rw1[19]
  PIN wd_in_rw1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 493.050 0.800 493.350 ;
    END
  END wd_in_rw1[20]
  PIN wd_in_rw1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 497.250 0.800 497.550 ;
    END
  END wd_in_rw1[21]
  PIN wd_in_rw1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 501.450 0.800 501.750 ;
    END
  END wd_in_rw1[22]
  PIN wd_in_rw1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 505.650 0.800 505.950 ;
    END
  END wd_in_rw1[23]
  PIN wd_in_rw1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 509.850 0.800 510.150 ;
    END
  END wd_in_rw1[24]
  PIN wd_in_rw1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 514.050 0.800 514.350 ;
    END
  END wd_in_rw1[25]
  PIN wd_in_rw1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 518.250 0.800 518.550 ;
    END
  END wd_in_rw1[26]
  PIN wd_in_rw1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 522.450 0.800 522.750 ;
    END
  END wd_in_rw1[27]
  PIN wd_in_rw1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 526.650 0.800 526.950 ;
    END
  END wd_in_rw1[28]
  PIN wd_in_rw1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 530.850 0.800 531.150 ;
    END
  END wd_in_rw1[29]
  PIN wd_in_rw1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 535.050 0.800 535.350 ;
    END
  END wd_in_rw1[30]
  PIN wd_in_rw1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 539.250 0.800 539.550 ;
    END
  END wd_in_rw1[31]
  PIN addr_rw1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 543.450 0.800 543.750 ;
    END
  END addr_rw1[0]
  PIN addr_rw1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 547.650 0.800 547.950 ;
    END
  END addr_rw1[1]
  PIN addr_rw1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 551.850 0.800 552.150 ;
    END
  END addr_rw1[2]
  PIN addr_rw1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 556.050 0.800 556.350 ;
    END
  END addr_rw1[3]
  PIN addr_rw1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 560.250 0.800 560.550 ;
    END
  END addr_rw1[4]
  PIN addr_rw1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 564.450 0.800 564.750 ;
    END
  END addr_rw1[5]
  PIN addr_rw1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 568.650 0.800 568.950 ;
    END
  END addr_rw1[6]
  PIN addr_rw1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 572.850 0.800 573.150 ;
    END
  END addr_rw1[7]
  PIN addr_rw1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 577.050 0.800 577.350 ;
    END
  END addr_rw1[8]
  PIN addr_r1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 581.250 0.800 581.550 ;
    END
  END addr_r1[0]
  PIN addr_r1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 585.450 0.800 585.750 ;
    END
  END addr_r1[1]
  PIN addr_r1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 589.650 0.800 589.950 ;
    END
  END addr_r1[2]
  PIN addr_r1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 593.850 0.800 594.150 ;
    END
  END addr_r1[3]
  PIN addr_r1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 598.050 0.800 598.350 ;
    END
  END addr_r1[4]
  PIN addr_r1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 602.250 0.800 602.550 ;
    END
  END addr_r1[5]
  PIN addr_r1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 606.450 0.800 606.750 ;
    END
  END addr_r1[6]
  PIN addr_r1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 610.650 0.800 610.950 ;
    END
  END addr_r1[7]
  PIN addr_r1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 614.850 0.800 615.150 ;
    END
  END addr_r1[8]
  PIN we_in_rw1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 619.050 0.800 619.350 ;
    END
  END we_in_rw1
  PIN ce_rw1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 623.250 0.800 623.550 ;
    END
  END ce_rw1
  PIN ce_r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 627.450 0.800 627.750 ;
    END
  END ce_r1
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 631.650 0.800 631.950 ;
    END
  END clk0
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 635.850 0.800 636.150 ;
    END
  END clk1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 5.400 6.000 6.600 538.000 ;
      RECT 15.000 6.000 16.200 538.000 ;
      RECT 24.600 6.000 25.800 538.000 ;
      RECT 34.200 6.000 35.400 538.000 ;
      RECT 43.800 6.000 45.000 538.000 ;
      RECT 53.400 6.000 54.600 538.000 ;
      RECT 63.000 6.000 64.200 538.000 ;
      RECT 72.600 6.000 73.800 538.000 ;
      RECT 82.200 6.000 83.400 538.000 ;
      RECT 91.800 6.000 93.000 538.000 ;
      RECT 101.400 6.000 102.600 538.000 ;
      RECT 111.000 6.000 112.200 538.000 ;
      RECT 120.600 6.000 121.800 538.000 ;
      RECT 130.200 6.000 131.400 538.000 ;
      RECT 139.800 6.000 141.000 538.000 ;
      RECT 149.400 6.000 150.600 538.000 ;
      RECT 159.000 6.000 160.200 538.000 ;
      RECT 168.600 6.000 169.800 538.000 ;
      RECT 178.200 6.000 179.400 538.000 ;
      RECT 187.800 6.000 189.000 538.000 ;
      RECT 197.400 6.000 198.600 538.000 ;
      RECT 207.000 6.000 208.200 538.000 ;
      RECT 216.600 6.000 217.800 538.000 ;
      RECT 226.200 6.000 227.400 538.000 ;
      RECT 235.800 6.000 237.000 538.000 ;
      RECT 245.400 6.000 246.600 538.000 ;
      RECT 255.000 6.000 256.200 538.000 ;
      RECT 264.600 6.000 265.800 538.000 ;
      RECT 274.200 6.000 275.400 538.000 ;
      RECT 283.800 6.000 285.000 538.000 ;
      RECT 293.400 6.000 294.600 538.000 ;
      RECT 303.000 6.000 304.200 538.000 ;
      RECT 312.600 6.000 313.800 538.000 ;
      RECT 322.200 6.000 323.400 538.000 ;
      RECT 331.800 6.000 333.000 538.000 ;
      RECT 341.400 6.000 342.600 538.000 ;
      RECT 351.000 6.000 352.200 538.000 ;
      RECT 360.600 6.000 361.800 538.000 ;
      RECT 370.200 6.000 371.400 538.000 ;
      RECT 379.800 6.000 381.000 538.000 ;
      RECT 389.400 6.000 390.600 538.000 ;
      RECT 399.000 6.000 400.200 538.000 ;
      RECT 408.600 6.000 409.800 538.000 ;
      RECT 418.200 6.000 419.400 538.000 ;
      RECT 427.800 6.000 429.000 538.000 ;
      RECT 437.400 6.000 438.600 538.000 ;
      RECT 447.000 6.000 448.200 538.000 ;
      RECT 456.600 6.000 457.800 538.000 ;
      RECT 466.200 6.000 467.400 538.000 ;
      RECT 475.800 6.000 477.000 538.000 ;
      RECT 485.400 6.000 486.600 538.000 ;
      RECT 495.000 6.000 496.200 538.000 ;
      RECT 504.600 6.000 505.800 538.000 ;
      RECT 514.200 6.000 515.400 538.000 ;
      RECT 523.800 6.000 525.000 538.000 ;
      RECT 533.400 6.000 534.600 538.000 ;
      RECT 543.000 6.000 544.200 538.000 ;
      RECT 552.600 6.000 553.800 538.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 10.200 6.000 11.400 538.000 ;
      RECT 19.800 6.000 21.000 538.000 ;
      RECT 29.400 6.000 30.600 538.000 ;
      RECT 39.000 6.000 40.200 538.000 ;
      RECT 48.600 6.000 49.800 538.000 ;
      RECT 58.200 6.000 59.400 538.000 ;
      RECT 67.800 6.000 69.000 538.000 ;
      RECT 77.400 6.000 78.600 538.000 ;
      RECT 87.000 6.000 88.200 538.000 ;
      RECT 96.600 6.000 97.800 538.000 ;
      RECT 106.200 6.000 107.400 538.000 ;
      RECT 115.800 6.000 117.000 538.000 ;
      RECT 125.400 6.000 126.600 538.000 ;
      RECT 135.000 6.000 136.200 538.000 ;
      RECT 144.600 6.000 145.800 538.000 ;
      RECT 154.200 6.000 155.400 538.000 ;
      RECT 163.800 6.000 165.000 538.000 ;
      RECT 173.400 6.000 174.600 538.000 ;
      RECT 183.000 6.000 184.200 538.000 ;
      RECT 192.600 6.000 193.800 538.000 ;
      RECT 202.200 6.000 203.400 538.000 ;
      RECT 211.800 6.000 213.000 538.000 ;
      RECT 221.400 6.000 222.600 538.000 ;
      RECT 231.000 6.000 232.200 538.000 ;
      RECT 240.600 6.000 241.800 538.000 ;
      RECT 250.200 6.000 251.400 538.000 ;
      RECT 259.800 6.000 261.000 538.000 ;
      RECT 269.400 6.000 270.600 538.000 ;
      RECT 279.000 6.000 280.200 538.000 ;
      RECT 288.600 6.000 289.800 538.000 ;
      RECT 298.200 6.000 299.400 538.000 ;
      RECT 307.800 6.000 309.000 538.000 ;
      RECT 317.400 6.000 318.600 538.000 ;
      RECT 327.000 6.000 328.200 538.000 ;
      RECT 336.600 6.000 337.800 538.000 ;
      RECT 346.200 6.000 347.400 538.000 ;
      RECT 355.800 6.000 357.000 538.000 ;
      RECT 365.400 6.000 366.600 538.000 ;
      RECT 375.000 6.000 376.200 538.000 ;
      RECT 384.600 6.000 385.800 538.000 ;
      RECT 394.200 6.000 395.400 538.000 ;
      RECT 403.800 6.000 405.000 538.000 ;
      RECT 413.400 6.000 414.600 538.000 ;
      RECT 423.000 6.000 424.200 538.000 ;
      RECT 432.600 6.000 433.800 538.000 ;
      RECT 442.200 6.000 443.400 538.000 ;
      RECT 451.800 6.000 453.000 538.000 ;
      RECT 461.400 6.000 462.600 538.000 ;
      RECT 471.000 6.000 472.200 538.000 ;
      RECT 480.600 6.000 481.800 538.000 ;
      RECT 490.200 6.000 491.400 538.000 ;
      RECT 499.800 6.000 501.000 538.000 ;
      RECT 509.400 6.000 510.600 538.000 ;
      RECT 519.000 6.000 520.200 538.000 ;
      RECT 528.600 6.000 529.800 538.000 ;
      RECT 538.200 6.000 539.400 538.000 ;
      RECT 547.800 6.000 549.000 538.000 ;
      RECT 557.400 6.000 558.600 538.000 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 568.100 544.000 ;
    LAYER met2 ;
    RECT 0 0 568.100 544.000 ;
    LAYER met3 ;
    RECT 0.800 0 568.100 544.000 ;
    RECT 0 0.000 0.800 5.850 ;
    RECT 0 6.150 0.800 10.050 ;
    RECT 0 10.350 0.800 14.250 ;
    RECT 0 14.550 0.800 18.450 ;
    RECT 0 18.750 0.800 22.650 ;
    RECT 0 22.950 0.800 26.850 ;
    RECT 0 27.150 0.800 31.050 ;
    RECT 0 31.350 0.800 35.250 ;
    RECT 0 35.550 0.800 39.450 ;
    RECT 0 39.750 0.800 43.650 ;
    RECT 0 43.950 0.800 47.850 ;
    RECT 0 48.150 0.800 52.050 ;
    RECT 0 52.350 0.800 56.250 ;
    RECT 0 56.550 0.800 60.450 ;
    RECT 0 60.750 0.800 64.650 ;
    RECT 0 64.950 0.800 68.850 ;
    RECT 0 69.150 0.800 73.050 ;
    RECT 0 73.350 0.800 77.250 ;
    RECT 0 77.550 0.800 81.450 ;
    RECT 0 81.750 0.800 85.650 ;
    RECT 0 85.950 0.800 89.850 ;
    RECT 0 90.150 0.800 94.050 ;
    RECT 0 94.350 0.800 98.250 ;
    RECT 0 98.550 0.800 102.450 ;
    RECT 0 102.750 0.800 106.650 ;
    RECT 0 106.950 0.800 110.850 ;
    RECT 0 111.150 0.800 115.050 ;
    RECT 0 115.350 0.800 119.250 ;
    RECT 0 119.550 0.800 123.450 ;
    RECT 0 123.750 0.800 127.650 ;
    RECT 0 127.950 0.800 131.850 ;
    RECT 0 132.150 0.800 136.050 ;
    RECT 0 136.350 0.800 140.250 ;
    RECT 0 140.550 0.800 144.450 ;
    RECT 0 144.750 0.800 148.650 ;
    RECT 0 148.950 0.800 152.850 ;
    RECT 0 153.150 0.800 157.050 ;
    RECT 0 157.350 0.800 161.250 ;
    RECT 0 161.550 0.800 165.450 ;
    RECT 0 165.750 0.800 169.650 ;
    RECT 0 169.950 0.800 173.850 ;
    RECT 0 174.150 0.800 178.050 ;
    RECT 0 178.350 0.800 182.250 ;
    RECT 0 182.550 0.800 186.450 ;
    RECT 0 186.750 0.800 190.650 ;
    RECT 0 190.950 0.800 194.850 ;
    RECT 0 195.150 0.800 199.050 ;
    RECT 0 199.350 0.800 203.250 ;
    RECT 0 203.550 0.800 207.450 ;
    RECT 0 207.750 0.800 211.650 ;
    RECT 0 211.950 0.800 215.850 ;
    RECT 0 216.150 0.800 220.050 ;
    RECT 0 220.350 0.800 224.250 ;
    RECT 0 224.550 0.800 228.450 ;
    RECT 0 228.750 0.800 232.650 ;
    RECT 0 232.950 0.800 236.850 ;
    RECT 0 237.150 0.800 241.050 ;
    RECT 0 241.350 0.800 245.250 ;
    RECT 0 245.550 0.800 249.450 ;
    RECT 0 249.750 0.800 253.650 ;
    RECT 0 253.950 0.800 257.850 ;
    RECT 0 258.150 0.800 262.050 ;
    RECT 0 262.350 0.800 266.250 ;
    RECT 0 266.550 0.800 270.450 ;
    RECT 0 270.750 0.800 274.650 ;
    RECT 0 274.950 0.800 278.850 ;
    RECT 0 279.150 0.800 283.050 ;
    RECT 0 283.350 0.800 287.250 ;
    RECT 0 287.550 0.800 291.450 ;
    RECT 0 291.750 0.800 295.650 ;
    RECT 0 295.950 0.800 299.850 ;
    RECT 0 300.150 0.800 304.050 ;
    RECT 0 304.350 0.800 308.250 ;
    RECT 0 308.550 0.800 312.450 ;
    RECT 0 312.750 0.800 316.650 ;
    RECT 0 316.950 0.800 320.850 ;
    RECT 0 321.150 0.800 325.050 ;
    RECT 0 325.350 0.800 329.250 ;
    RECT 0 329.550 0.800 333.450 ;
    RECT 0 333.750 0.800 337.650 ;
    RECT 0 337.950 0.800 341.850 ;
    RECT 0 342.150 0.800 346.050 ;
    RECT 0 346.350 0.800 350.250 ;
    RECT 0 350.550 0.800 354.450 ;
    RECT 0 354.750 0.800 358.650 ;
    RECT 0 358.950 0.800 362.850 ;
    RECT 0 363.150 0.800 367.050 ;
    RECT 0 367.350 0.800 371.250 ;
    RECT 0 371.550 0.800 375.450 ;
    RECT 0 375.750 0.800 379.650 ;
    RECT 0 379.950 0.800 383.850 ;
    RECT 0 384.150 0.800 388.050 ;
    RECT 0 388.350 0.800 392.250 ;
    RECT 0 392.550 0.800 396.450 ;
    RECT 0 396.750 0.800 400.650 ;
    RECT 0 400.950 0.800 404.850 ;
    RECT 0 405.150 0.800 409.050 ;
    RECT 0 409.350 0.800 413.250 ;
    RECT 0 413.550 0.800 417.450 ;
    RECT 0 417.750 0.800 421.650 ;
    RECT 0 421.950 0.800 425.850 ;
    RECT 0 426.150 0.800 430.050 ;
    RECT 0 430.350 0.800 434.250 ;
    RECT 0 434.550 0.800 438.450 ;
    RECT 0 438.750 0.800 442.650 ;
    RECT 0 442.950 0.800 446.850 ;
    RECT 0 447.150 0.800 451.050 ;
    RECT 0 451.350 0.800 455.250 ;
    RECT 0 455.550 0.800 544.000 ;
    LAYER met4 ;
    RECT 0 0 568.100 6.000 ;
    RECT 0 538.000 568.100 544.000 ;
    RECT 0.000 6.000 5.400 538.000 ;
    RECT 6.600 6.000 10.200 538.000 ;
    RECT 11.400 6.000 15.000 538.000 ;
    RECT 16.200 6.000 19.800 538.000 ;
    RECT 21.000 6.000 24.600 538.000 ;
    RECT 25.800 6.000 29.400 538.000 ;
    RECT 30.600 6.000 34.200 538.000 ;
    RECT 35.400 6.000 39.000 538.000 ;
    RECT 40.200 6.000 43.800 538.000 ;
    RECT 45.000 6.000 48.600 538.000 ;
    RECT 49.800 6.000 53.400 538.000 ;
    RECT 54.600 6.000 58.200 538.000 ;
    RECT 59.400 6.000 63.000 538.000 ;
    RECT 64.200 6.000 67.800 538.000 ;
    RECT 69.000 6.000 72.600 538.000 ;
    RECT 73.800 6.000 77.400 538.000 ;
    RECT 78.600 6.000 82.200 538.000 ;
    RECT 83.400 6.000 87.000 538.000 ;
    RECT 88.200 6.000 91.800 538.000 ;
    RECT 93.000 6.000 96.600 538.000 ;
    RECT 97.800 6.000 101.400 538.000 ;
    RECT 102.600 6.000 106.200 538.000 ;
    RECT 107.400 6.000 111.000 538.000 ;
    RECT 112.200 6.000 115.800 538.000 ;
    RECT 117.000 6.000 120.600 538.000 ;
    RECT 121.800 6.000 125.400 538.000 ;
    RECT 126.600 6.000 130.200 538.000 ;
    RECT 131.400 6.000 135.000 538.000 ;
    RECT 136.200 6.000 139.800 538.000 ;
    RECT 141.000 6.000 144.600 538.000 ;
    RECT 145.800 6.000 149.400 538.000 ;
    RECT 150.600 6.000 154.200 538.000 ;
    RECT 155.400 6.000 159.000 538.000 ;
    RECT 160.200 6.000 163.800 538.000 ;
    RECT 165.000 6.000 168.600 538.000 ;
    RECT 169.800 6.000 173.400 538.000 ;
    RECT 174.600 6.000 178.200 538.000 ;
    RECT 179.400 6.000 183.000 538.000 ;
    RECT 184.200 6.000 187.800 538.000 ;
    RECT 189.000 6.000 192.600 538.000 ;
    RECT 193.800 6.000 197.400 538.000 ;
    RECT 198.600 6.000 202.200 538.000 ;
    RECT 203.400 6.000 207.000 538.000 ;
    RECT 208.200 6.000 211.800 538.000 ;
    RECT 213.000 6.000 216.600 538.000 ;
    RECT 217.800 6.000 221.400 538.000 ;
    RECT 222.600 6.000 226.200 538.000 ;
    RECT 227.400 6.000 231.000 538.000 ;
    RECT 232.200 6.000 235.800 538.000 ;
    RECT 237.000 6.000 240.600 538.000 ;
    RECT 241.800 6.000 245.400 538.000 ;
    RECT 246.600 6.000 250.200 538.000 ;
    RECT 251.400 6.000 255.000 538.000 ;
    RECT 256.200 6.000 259.800 538.000 ;
    RECT 261.000 6.000 264.600 538.000 ;
    RECT 265.800 6.000 269.400 538.000 ;
    RECT 270.600 6.000 274.200 538.000 ;
    RECT 275.400 6.000 279.000 538.000 ;
    RECT 280.200 6.000 283.800 538.000 ;
    RECT 285.000 6.000 288.600 538.000 ;
    RECT 289.800 6.000 293.400 538.000 ;
    RECT 294.600 6.000 298.200 538.000 ;
    RECT 299.400 6.000 303.000 538.000 ;
    RECT 304.200 6.000 307.800 538.000 ;
    RECT 309.000 6.000 312.600 538.000 ;
    RECT 313.800 6.000 317.400 538.000 ;
    RECT 318.600 6.000 322.200 538.000 ;
    RECT 323.400 6.000 327.000 538.000 ;
    RECT 328.200 6.000 331.800 538.000 ;
    RECT 333.000 6.000 336.600 538.000 ;
    RECT 337.800 6.000 341.400 538.000 ;
    RECT 342.600 6.000 346.200 538.000 ;
    RECT 347.400 6.000 351.000 538.000 ;
    RECT 352.200 6.000 355.800 538.000 ;
    RECT 357.000 6.000 360.600 538.000 ;
    RECT 361.800 6.000 365.400 538.000 ;
    RECT 366.600 6.000 370.200 538.000 ;
    RECT 371.400 6.000 375.000 538.000 ;
    RECT 376.200 6.000 379.800 538.000 ;
    RECT 381.000 6.000 384.600 538.000 ;
    RECT 385.800 6.000 389.400 538.000 ;
    RECT 390.600 6.000 394.200 538.000 ;
    RECT 395.400 6.000 399.000 538.000 ;
    RECT 400.200 6.000 403.800 538.000 ;
    RECT 405.000 6.000 408.600 538.000 ;
    RECT 409.800 6.000 413.400 538.000 ;
    RECT 414.600 6.000 418.200 538.000 ;
    RECT 419.400 6.000 423.000 538.000 ;
    RECT 424.200 6.000 427.800 538.000 ;
    RECT 429.000 6.000 432.600 538.000 ;
    RECT 433.800 6.000 437.400 538.000 ;
    RECT 438.600 6.000 442.200 538.000 ;
    RECT 443.400 6.000 447.000 538.000 ;
    RECT 448.200 6.000 451.800 538.000 ;
    RECT 453.000 6.000 456.600 538.000 ;
    RECT 457.800 6.000 461.400 538.000 ;
    RECT 462.600 6.000 466.200 538.000 ;
    RECT 467.400 6.000 471.000 538.000 ;
    RECT 472.200 6.000 475.800 538.000 ;
    RECT 477.000 6.000 480.600 538.000 ;
    RECT 481.800 6.000 485.400 538.000 ;
    RECT 486.600 6.000 490.200 538.000 ;
    RECT 491.400 6.000 495.000 538.000 ;
    RECT 496.200 6.000 499.800 538.000 ;
    RECT 501.000 6.000 504.600 538.000 ;
    RECT 505.800 6.000 509.400 538.000 ;
    RECT 510.600 6.000 514.200 538.000 ;
    RECT 515.400 6.000 519.000 538.000 ;
    RECT 520.200 6.000 523.800 538.000 ;
    RECT 525.000 6.000 528.600 538.000 ;
    RECT 529.800 6.000 533.400 538.000 ;
    RECT 534.600 6.000 538.200 538.000 ;
    RECT 539.400 6.000 543.000 538.000 ;
    RECT 544.200 6.000 547.800 538.000 ;
    RECT 549.000 6.000 552.600 538.000 ;
    RECT 553.800 6.000 557.400 538.000 ;
    RECT 558.600 6.000 568.100 538.000 ;
    LAYER OVERLAP ;
    RECT 0 0 568.100 544.000 ;
  END
END liteeth_1rw1r_32w384d_32_sram

END LIBRARY
