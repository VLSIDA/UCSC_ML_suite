VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_512x256_1r1w
  FOREIGN fakeram_512x256_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 689.130 BY 767.200 ;
  CLASS BLOCK ;
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 0.805 0.140 0.875 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.405 0.140 6.475 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.005 0.140 12.075 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.140 17.675 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.205 0.140 23.275 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.805 0.140 28.875 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.140 34.475 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.005 0.140 40.075 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.605 0.140 45.675 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.140 51.275 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.805 0.140 56.875 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.405 0.140 62.475 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.005 0.140 68.075 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.605 0.140 73.675 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.205 0.140 79.275 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.140 84.875 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.405 0.140 90.475 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.005 0.140 96.075 ;
    END
  END w0_wd_in[17]
  PIN w0_wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.605 0.140 101.675 ;
    END
  END w0_wd_in[18]
  PIN w0_wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.205 0.140 107.275 ;
    END
  END w0_wd_in[19]
  PIN w0_wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.805 0.140 112.875 ;
    END
  END w0_wd_in[20]
  PIN w0_wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.405 0.140 118.475 ;
    END
  END w0_wd_in[21]
  PIN w0_wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.005 0.140 124.075 ;
    END
  END w0_wd_in[22]
  PIN w0_wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.605 0.140 129.675 ;
    END
  END w0_wd_in[23]
  PIN w0_wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.205 0.140 135.275 ;
    END
  END w0_wd_in[24]
  PIN w0_wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.805 0.140 140.875 ;
    END
  END w0_wd_in[25]
  PIN w0_wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.405 0.140 146.475 ;
    END
  END w0_wd_in[26]
  PIN w0_wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.005 0.140 152.075 ;
    END
  END w0_wd_in[27]
  PIN w0_wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.605 0.140 157.675 ;
    END
  END w0_wd_in[28]
  PIN w0_wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.205 0.140 163.275 ;
    END
  END w0_wd_in[29]
  PIN w0_wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.805 0.140 168.875 ;
    END
  END w0_wd_in[30]
  PIN w0_wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.405 0.140 174.475 ;
    END
  END w0_wd_in[31]
  PIN w0_wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.005 0.140 180.075 ;
    END
  END w0_wd_in[32]
  PIN w0_wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.605 0.140 185.675 ;
    END
  END w0_wd_in[33]
  PIN w0_wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.205 0.140 191.275 ;
    END
  END w0_wd_in[34]
  PIN w0_wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.805 0.140 196.875 ;
    END
  END w0_wd_in[35]
  PIN w0_wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.405 0.140 202.475 ;
    END
  END w0_wd_in[36]
  PIN w0_wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.005 0.140 208.075 ;
    END
  END w0_wd_in[37]
  PIN w0_wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.605 0.140 213.675 ;
    END
  END w0_wd_in[38]
  PIN w0_wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.205 0.140 219.275 ;
    END
  END w0_wd_in[39]
  PIN w0_wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.805 0.140 224.875 ;
    END
  END w0_wd_in[40]
  PIN w0_wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.405 0.140 230.475 ;
    END
  END w0_wd_in[41]
  PIN w0_wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.005 0.140 236.075 ;
    END
  END w0_wd_in[42]
  PIN w0_wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.605 0.140 241.675 ;
    END
  END w0_wd_in[43]
  PIN w0_wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.205 0.140 247.275 ;
    END
  END w0_wd_in[44]
  PIN w0_wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.805 0.140 252.875 ;
    END
  END w0_wd_in[45]
  PIN w0_wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.405 0.140 258.475 ;
    END
  END w0_wd_in[46]
  PIN w0_wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.005 0.140 264.075 ;
    END
  END w0_wd_in[47]
  PIN w0_wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.605 0.140 269.675 ;
    END
  END w0_wd_in[48]
  PIN w0_wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.205 0.140 275.275 ;
    END
  END w0_wd_in[49]
  PIN w0_wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.805 0.140 280.875 ;
    END
  END w0_wd_in[50]
  PIN w0_wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.405 0.140 286.475 ;
    END
  END w0_wd_in[51]
  PIN w0_wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.005 0.140 292.075 ;
    END
  END w0_wd_in[52]
  PIN w0_wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.605 0.140 297.675 ;
    END
  END w0_wd_in[53]
  PIN w0_wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.205 0.140 303.275 ;
    END
  END w0_wd_in[54]
  PIN w0_wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.805 0.140 308.875 ;
    END
  END w0_wd_in[55]
  PIN w0_wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.405 0.140 314.475 ;
    END
  END w0_wd_in[56]
  PIN w0_wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.005 0.140 320.075 ;
    END
  END w0_wd_in[57]
  PIN w0_wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.605 0.140 325.675 ;
    END
  END w0_wd_in[58]
  PIN w0_wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.205 0.140 331.275 ;
    END
  END w0_wd_in[59]
  PIN w0_wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.805 0.140 336.875 ;
    END
  END w0_wd_in[60]
  PIN w0_wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.405 0.140 342.475 ;
    END
  END w0_wd_in[61]
  PIN w0_wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.005 0.140 348.075 ;
    END
  END w0_wd_in[62]
  PIN w0_wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.605 0.140 353.675 ;
    END
  END w0_wd_in[63]
  PIN w0_wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.205 0.140 359.275 ;
    END
  END w0_wd_in[64]
  PIN w0_wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.805 0.140 364.875 ;
    END
  END w0_wd_in[65]
  PIN w0_wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.405 0.140 370.475 ;
    END
  END w0_wd_in[66]
  PIN w0_wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.005 0.140 376.075 ;
    END
  END w0_wd_in[67]
  PIN w0_wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.605 0.140 381.675 ;
    END
  END w0_wd_in[68]
  PIN w0_wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.205 0.140 387.275 ;
    END
  END w0_wd_in[69]
  PIN w0_wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.805 0.140 392.875 ;
    END
  END w0_wd_in[70]
  PIN w0_wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.405 0.140 398.475 ;
    END
  END w0_wd_in[71]
  PIN w0_wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 404.005 0.140 404.075 ;
    END
  END w0_wd_in[72]
  PIN w0_wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 409.605 0.140 409.675 ;
    END
  END w0_wd_in[73]
  PIN w0_wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 415.205 0.140 415.275 ;
    END
  END w0_wd_in[74]
  PIN w0_wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 420.805 0.140 420.875 ;
    END
  END w0_wd_in[75]
  PIN w0_wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 426.405 0.140 426.475 ;
    END
  END w0_wd_in[76]
  PIN w0_wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 432.005 0.140 432.075 ;
    END
  END w0_wd_in[77]
  PIN w0_wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 437.605 0.140 437.675 ;
    END
  END w0_wd_in[78]
  PIN w0_wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 443.205 0.140 443.275 ;
    END
  END w0_wd_in[79]
  PIN w0_wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 448.805 0.140 448.875 ;
    END
  END w0_wd_in[80]
  PIN w0_wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 454.405 0.140 454.475 ;
    END
  END w0_wd_in[81]
  PIN w0_wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 460.005 0.140 460.075 ;
    END
  END w0_wd_in[82]
  PIN w0_wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 465.605 0.140 465.675 ;
    END
  END w0_wd_in[83]
  PIN w0_wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 471.205 0.140 471.275 ;
    END
  END w0_wd_in[84]
  PIN w0_wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 476.805 0.140 476.875 ;
    END
  END w0_wd_in[85]
  PIN w0_wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 482.405 0.140 482.475 ;
    END
  END w0_wd_in[86]
  PIN w0_wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 488.005 0.140 488.075 ;
    END
  END w0_wd_in[87]
  PIN w0_wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 493.605 0.140 493.675 ;
    END
  END w0_wd_in[88]
  PIN w0_wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 499.205 0.140 499.275 ;
    END
  END w0_wd_in[89]
  PIN w0_wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 504.805 0.140 504.875 ;
    END
  END w0_wd_in[90]
  PIN w0_wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.405 0.140 510.475 ;
    END
  END w0_wd_in[91]
  PIN w0_wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.005 0.140 516.075 ;
    END
  END w0_wd_in[92]
  PIN w0_wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.605 0.140 521.675 ;
    END
  END w0_wd_in[93]
  PIN w0_wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.205 0.140 527.275 ;
    END
  END w0_wd_in[94]
  PIN w0_wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.805 0.140 532.875 ;
    END
  END w0_wd_in[95]
  PIN w0_wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.405 0.140 538.475 ;
    END
  END w0_wd_in[96]
  PIN w0_wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.005 0.140 544.075 ;
    END
  END w0_wd_in[97]
  PIN w0_wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.605 0.140 549.675 ;
    END
  END w0_wd_in[98]
  PIN w0_wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.205 0.140 555.275 ;
    END
  END w0_wd_in[99]
  PIN w0_wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.805 0.140 560.875 ;
    END
  END w0_wd_in[100]
  PIN w0_wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.405 0.140 566.475 ;
    END
  END w0_wd_in[101]
  PIN w0_wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.005 0.140 572.075 ;
    END
  END w0_wd_in[102]
  PIN w0_wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.605 0.140 577.675 ;
    END
  END w0_wd_in[103]
  PIN w0_wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.205 0.140 583.275 ;
    END
  END w0_wd_in[104]
  PIN w0_wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.805 0.140 588.875 ;
    END
  END w0_wd_in[105]
  PIN w0_wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.405 0.140 594.475 ;
    END
  END w0_wd_in[106]
  PIN w0_wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.005 0.140 600.075 ;
    END
  END w0_wd_in[107]
  PIN w0_wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.605 0.140 605.675 ;
    END
  END w0_wd_in[108]
  PIN w0_wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.205 0.140 611.275 ;
    END
  END w0_wd_in[109]
  PIN w0_wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.805 0.140 616.875 ;
    END
  END w0_wd_in[110]
  PIN w0_wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.405 0.140 622.475 ;
    END
  END w0_wd_in[111]
  PIN w0_wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.005 0.140 628.075 ;
    END
  END w0_wd_in[112]
  PIN w0_wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.605 0.140 633.675 ;
    END
  END w0_wd_in[113]
  PIN w0_wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 639.205 0.140 639.275 ;
    END
  END w0_wd_in[114]
  PIN w0_wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 644.805 0.140 644.875 ;
    END
  END w0_wd_in[115]
  PIN w0_wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 650.405 0.140 650.475 ;
    END
  END w0_wd_in[116]
  PIN w0_wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.005 0.140 656.075 ;
    END
  END w0_wd_in[117]
  PIN w0_wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.605 0.140 661.675 ;
    END
  END w0_wd_in[118]
  PIN w0_wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.205 0.140 667.275 ;
    END
  END w0_wd_in[119]
  PIN w0_wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.805 0.140 672.875 ;
    END
  END w0_wd_in[120]
  PIN w0_wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.405 0.140 678.475 ;
    END
  END w0_wd_in[121]
  PIN w0_wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.005 0.140 684.075 ;
    END
  END w0_wd_in[122]
  PIN w0_wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.605 0.140 689.675 ;
    END
  END w0_wd_in[123]
  PIN w0_wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 695.205 0.140 695.275 ;
    END
  END w0_wd_in[124]
  PIN w0_wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 700.805 0.140 700.875 ;
    END
  END w0_wd_in[125]
  PIN w0_wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.405 0.140 706.475 ;
    END
  END w0_wd_in[126]
  PIN w0_wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.005 0.140 712.075 ;
    END
  END w0_wd_in[127]
  PIN w0_wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 0.805 689.130 0.875 ;
    END
  END w0_wd_in[128]
  PIN w0_wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 6.405 689.130 6.475 ;
    END
  END w0_wd_in[129]
  PIN w0_wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 12.005 689.130 12.075 ;
    END
  END w0_wd_in[130]
  PIN w0_wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 17.605 689.130 17.675 ;
    END
  END w0_wd_in[131]
  PIN w0_wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 23.205 689.130 23.275 ;
    END
  END w0_wd_in[132]
  PIN w0_wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 28.805 689.130 28.875 ;
    END
  END w0_wd_in[133]
  PIN w0_wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 34.405 689.130 34.475 ;
    END
  END w0_wd_in[134]
  PIN w0_wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 40.005 689.130 40.075 ;
    END
  END w0_wd_in[135]
  PIN w0_wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 45.605 689.130 45.675 ;
    END
  END w0_wd_in[136]
  PIN w0_wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 51.205 689.130 51.275 ;
    END
  END w0_wd_in[137]
  PIN w0_wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 56.805 689.130 56.875 ;
    END
  END w0_wd_in[138]
  PIN w0_wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 62.405 689.130 62.475 ;
    END
  END w0_wd_in[139]
  PIN w0_wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 68.005 689.130 68.075 ;
    END
  END w0_wd_in[140]
  PIN w0_wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 73.605 689.130 73.675 ;
    END
  END w0_wd_in[141]
  PIN w0_wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 79.205 689.130 79.275 ;
    END
  END w0_wd_in[142]
  PIN w0_wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 84.805 689.130 84.875 ;
    END
  END w0_wd_in[143]
  PIN w0_wd_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 90.405 689.130 90.475 ;
    END
  END w0_wd_in[144]
  PIN w0_wd_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 96.005 689.130 96.075 ;
    END
  END w0_wd_in[145]
  PIN w0_wd_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 101.605 689.130 101.675 ;
    END
  END w0_wd_in[146]
  PIN w0_wd_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 107.205 689.130 107.275 ;
    END
  END w0_wd_in[147]
  PIN w0_wd_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 112.805 689.130 112.875 ;
    END
  END w0_wd_in[148]
  PIN w0_wd_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 118.405 689.130 118.475 ;
    END
  END w0_wd_in[149]
  PIN w0_wd_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 124.005 689.130 124.075 ;
    END
  END w0_wd_in[150]
  PIN w0_wd_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 129.605 689.130 129.675 ;
    END
  END w0_wd_in[151]
  PIN w0_wd_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 135.205 689.130 135.275 ;
    END
  END w0_wd_in[152]
  PIN w0_wd_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 140.805 689.130 140.875 ;
    END
  END w0_wd_in[153]
  PIN w0_wd_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 146.405 689.130 146.475 ;
    END
  END w0_wd_in[154]
  PIN w0_wd_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 152.005 689.130 152.075 ;
    END
  END w0_wd_in[155]
  PIN w0_wd_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 157.605 689.130 157.675 ;
    END
  END w0_wd_in[156]
  PIN w0_wd_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 163.205 689.130 163.275 ;
    END
  END w0_wd_in[157]
  PIN w0_wd_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 168.805 689.130 168.875 ;
    END
  END w0_wd_in[158]
  PIN w0_wd_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 174.405 689.130 174.475 ;
    END
  END w0_wd_in[159]
  PIN w0_wd_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 180.005 689.130 180.075 ;
    END
  END w0_wd_in[160]
  PIN w0_wd_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 185.605 689.130 185.675 ;
    END
  END w0_wd_in[161]
  PIN w0_wd_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 191.205 689.130 191.275 ;
    END
  END w0_wd_in[162]
  PIN w0_wd_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 196.805 689.130 196.875 ;
    END
  END w0_wd_in[163]
  PIN w0_wd_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 202.405 689.130 202.475 ;
    END
  END w0_wd_in[164]
  PIN w0_wd_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 208.005 689.130 208.075 ;
    END
  END w0_wd_in[165]
  PIN w0_wd_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 213.605 689.130 213.675 ;
    END
  END w0_wd_in[166]
  PIN w0_wd_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 219.205 689.130 219.275 ;
    END
  END w0_wd_in[167]
  PIN w0_wd_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 224.805 689.130 224.875 ;
    END
  END w0_wd_in[168]
  PIN w0_wd_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 230.405 689.130 230.475 ;
    END
  END w0_wd_in[169]
  PIN w0_wd_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 236.005 689.130 236.075 ;
    END
  END w0_wd_in[170]
  PIN w0_wd_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 241.605 689.130 241.675 ;
    END
  END w0_wd_in[171]
  PIN w0_wd_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 247.205 689.130 247.275 ;
    END
  END w0_wd_in[172]
  PIN w0_wd_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 252.805 689.130 252.875 ;
    END
  END w0_wd_in[173]
  PIN w0_wd_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 258.405 689.130 258.475 ;
    END
  END w0_wd_in[174]
  PIN w0_wd_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 264.005 689.130 264.075 ;
    END
  END w0_wd_in[175]
  PIN w0_wd_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 269.605 689.130 269.675 ;
    END
  END w0_wd_in[176]
  PIN w0_wd_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 275.205 689.130 275.275 ;
    END
  END w0_wd_in[177]
  PIN w0_wd_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 280.805 689.130 280.875 ;
    END
  END w0_wd_in[178]
  PIN w0_wd_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 286.405 689.130 286.475 ;
    END
  END w0_wd_in[179]
  PIN w0_wd_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 292.005 689.130 292.075 ;
    END
  END w0_wd_in[180]
  PIN w0_wd_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 297.605 689.130 297.675 ;
    END
  END w0_wd_in[181]
  PIN w0_wd_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 303.205 689.130 303.275 ;
    END
  END w0_wd_in[182]
  PIN w0_wd_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 308.805 689.130 308.875 ;
    END
  END w0_wd_in[183]
  PIN w0_wd_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 314.405 689.130 314.475 ;
    END
  END w0_wd_in[184]
  PIN w0_wd_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 320.005 689.130 320.075 ;
    END
  END w0_wd_in[185]
  PIN w0_wd_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 325.605 689.130 325.675 ;
    END
  END w0_wd_in[186]
  PIN w0_wd_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 331.205 689.130 331.275 ;
    END
  END w0_wd_in[187]
  PIN w0_wd_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 336.805 689.130 336.875 ;
    END
  END w0_wd_in[188]
  PIN w0_wd_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 342.405 689.130 342.475 ;
    END
  END w0_wd_in[189]
  PIN w0_wd_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 348.005 689.130 348.075 ;
    END
  END w0_wd_in[190]
  PIN w0_wd_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 353.605 689.130 353.675 ;
    END
  END w0_wd_in[191]
  PIN w0_wd_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 359.205 689.130 359.275 ;
    END
  END w0_wd_in[192]
  PIN w0_wd_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 364.805 689.130 364.875 ;
    END
  END w0_wd_in[193]
  PIN w0_wd_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 370.405 689.130 370.475 ;
    END
  END w0_wd_in[194]
  PIN w0_wd_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 376.005 689.130 376.075 ;
    END
  END w0_wd_in[195]
  PIN w0_wd_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 381.605 689.130 381.675 ;
    END
  END w0_wd_in[196]
  PIN w0_wd_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 387.205 689.130 387.275 ;
    END
  END w0_wd_in[197]
  PIN w0_wd_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 392.805 689.130 392.875 ;
    END
  END w0_wd_in[198]
  PIN w0_wd_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 398.405 689.130 398.475 ;
    END
  END w0_wd_in[199]
  PIN w0_wd_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 404.005 689.130 404.075 ;
    END
  END w0_wd_in[200]
  PIN w0_wd_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 409.605 689.130 409.675 ;
    END
  END w0_wd_in[201]
  PIN w0_wd_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 415.205 689.130 415.275 ;
    END
  END w0_wd_in[202]
  PIN w0_wd_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 420.805 689.130 420.875 ;
    END
  END w0_wd_in[203]
  PIN w0_wd_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 426.405 689.130 426.475 ;
    END
  END w0_wd_in[204]
  PIN w0_wd_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 432.005 689.130 432.075 ;
    END
  END w0_wd_in[205]
  PIN w0_wd_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 437.605 689.130 437.675 ;
    END
  END w0_wd_in[206]
  PIN w0_wd_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 443.205 689.130 443.275 ;
    END
  END w0_wd_in[207]
  PIN w0_wd_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 448.805 689.130 448.875 ;
    END
  END w0_wd_in[208]
  PIN w0_wd_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 454.405 689.130 454.475 ;
    END
  END w0_wd_in[209]
  PIN w0_wd_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 460.005 689.130 460.075 ;
    END
  END w0_wd_in[210]
  PIN w0_wd_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 465.605 689.130 465.675 ;
    END
  END w0_wd_in[211]
  PIN w0_wd_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 471.205 689.130 471.275 ;
    END
  END w0_wd_in[212]
  PIN w0_wd_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 476.805 689.130 476.875 ;
    END
  END w0_wd_in[213]
  PIN w0_wd_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 482.405 689.130 482.475 ;
    END
  END w0_wd_in[214]
  PIN w0_wd_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 488.005 689.130 488.075 ;
    END
  END w0_wd_in[215]
  PIN w0_wd_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 493.605 689.130 493.675 ;
    END
  END w0_wd_in[216]
  PIN w0_wd_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 499.205 689.130 499.275 ;
    END
  END w0_wd_in[217]
  PIN w0_wd_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 504.805 689.130 504.875 ;
    END
  END w0_wd_in[218]
  PIN w0_wd_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 510.405 689.130 510.475 ;
    END
  END w0_wd_in[219]
  PIN w0_wd_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 516.005 689.130 516.075 ;
    END
  END w0_wd_in[220]
  PIN w0_wd_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 521.605 689.130 521.675 ;
    END
  END w0_wd_in[221]
  PIN w0_wd_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 527.205 689.130 527.275 ;
    END
  END w0_wd_in[222]
  PIN w0_wd_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 532.805 689.130 532.875 ;
    END
  END w0_wd_in[223]
  PIN w0_wd_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 538.405 689.130 538.475 ;
    END
  END w0_wd_in[224]
  PIN w0_wd_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 544.005 689.130 544.075 ;
    END
  END w0_wd_in[225]
  PIN w0_wd_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 549.605 689.130 549.675 ;
    END
  END w0_wd_in[226]
  PIN w0_wd_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 555.205 689.130 555.275 ;
    END
  END w0_wd_in[227]
  PIN w0_wd_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 560.805 689.130 560.875 ;
    END
  END w0_wd_in[228]
  PIN w0_wd_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 566.405 689.130 566.475 ;
    END
  END w0_wd_in[229]
  PIN w0_wd_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 572.005 689.130 572.075 ;
    END
  END w0_wd_in[230]
  PIN w0_wd_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 577.605 689.130 577.675 ;
    END
  END w0_wd_in[231]
  PIN w0_wd_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 583.205 689.130 583.275 ;
    END
  END w0_wd_in[232]
  PIN w0_wd_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 588.805 689.130 588.875 ;
    END
  END w0_wd_in[233]
  PIN w0_wd_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 594.405 689.130 594.475 ;
    END
  END w0_wd_in[234]
  PIN w0_wd_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 600.005 689.130 600.075 ;
    END
  END w0_wd_in[235]
  PIN w0_wd_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 605.605 689.130 605.675 ;
    END
  END w0_wd_in[236]
  PIN w0_wd_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 611.205 689.130 611.275 ;
    END
  END w0_wd_in[237]
  PIN w0_wd_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 616.805 689.130 616.875 ;
    END
  END w0_wd_in[238]
  PIN w0_wd_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 622.405 689.130 622.475 ;
    END
  END w0_wd_in[239]
  PIN w0_wd_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 628.005 689.130 628.075 ;
    END
  END w0_wd_in[240]
  PIN w0_wd_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 633.605 689.130 633.675 ;
    END
  END w0_wd_in[241]
  PIN w0_wd_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 639.205 689.130 639.275 ;
    END
  END w0_wd_in[242]
  PIN w0_wd_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 644.805 689.130 644.875 ;
    END
  END w0_wd_in[243]
  PIN w0_wd_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 650.405 689.130 650.475 ;
    END
  END w0_wd_in[244]
  PIN w0_wd_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 656.005 689.130 656.075 ;
    END
  END w0_wd_in[245]
  PIN w0_wd_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 661.605 689.130 661.675 ;
    END
  END w0_wd_in[246]
  PIN w0_wd_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 667.205 689.130 667.275 ;
    END
  END w0_wd_in[247]
  PIN w0_wd_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 672.805 689.130 672.875 ;
    END
  END w0_wd_in[248]
  PIN w0_wd_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 678.405 689.130 678.475 ;
    END
  END w0_wd_in[249]
  PIN w0_wd_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 684.005 689.130 684.075 ;
    END
  END w0_wd_in[250]
  PIN w0_wd_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 689.605 689.130 689.675 ;
    END
  END w0_wd_in[251]
  PIN w0_wd_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 695.205 689.130 695.275 ;
    END
  END w0_wd_in[252]
  PIN w0_wd_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 700.805 689.130 700.875 ;
    END
  END w0_wd_in[253]
  PIN w0_wd_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 706.405 689.130 706.475 ;
    END
  END w0_wd_in[254]
  PIN w0_wd_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 712.005 689.130 712.075 ;
    END
  END w0_wd_in[255]
  PIN w0_wd_in[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1.105 0.000 1.175 0.140 ;
    END
  END w0_wd_in[256]
  PIN w0_wd_in[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 2.435 0.000 2.505 0.140 ;
    END
  END w0_wd_in[257]
  PIN w0_wd_in[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 3.765 0.000 3.835 0.140 ;
    END
  END w0_wd_in[258]
  PIN w0_wd_in[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 5.095 0.000 5.165 0.140 ;
    END
  END w0_wd_in[259]
  PIN w0_wd_in[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 6.425 0.000 6.495 0.140 ;
    END
  END w0_wd_in[260]
  PIN w0_wd_in[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 7.755 0.000 7.825 0.140 ;
    END
  END w0_wd_in[261]
  PIN w0_wd_in[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 9.085 0.000 9.155 0.140 ;
    END
  END w0_wd_in[262]
  PIN w0_wd_in[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 10.415 0.000 10.485 0.140 ;
    END
  END w0_wd_in[263]
  PIN w0_wd_in[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 11.745 0.000 11.815 0.140 ;
    END
  END w0_wd_in[264]
  PIN w0_wd_in[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 13.075 0.000 13.145 0.140 ;
    END
  END w0_wd_in[265]
  PIN w0_wd_in[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 14.405 0.000 14.475 0.140 ;
    END
  END w0_wd_in[266]
  PIN w0_wd_in[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 15.735 0.000 15.805 0.140 ;
    END
  END w0_wd_in[267]
  PIN w0_wd_in[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 17.065 0.000 17.135 0.140 ;
    END
  END w0_wd_in[268]
  PIN w0_wd_in[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 18.395 0.000 18.465 0.140 ;
    END
  END w0_wd_in[269]
  PIN w0_wd_in[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 19.725 0.000 19.795 0.140 ;
    END
  END w0_wd_in[270]
  PIN w0_wd_in[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 21.055 0.000 21.125 0.140 ;
    END
  END w0_wd_in[271]
  PIN w0_wd_in[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 22.385 0.000 22.455 0.140 ;
    END
  END w0_wd_in[272]
  PIN w0_wd_in[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 23.715 0.000 23.785 0.140 ;
    END
  END w0_wd_in[273]
  PIN w0_wd_in[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 25.045 0.000 25.115 0.140 ;
    END
  END w0_wd_in[274]
  PIN w0_wd_in[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 26.375 0.000 26.445 0.140 ;
    END
  END w0_wd_in[275]
  PIN w0_wd_in[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 27.705 0.000 27.775 0.140 ;
    END
  END w0_wd_in[276]
  PIN w0_wd_in[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 29.035 0.000 29.105 0.140 ;
    END
  END w0_wd_in[277]
  PIN w0_wd_in[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 30.365 0.000 30.435 0.140 ;
    END
  END w0_wd_in[278]
  PIN w0_wd_in[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 31.695 0.000 31.765 0.140 ;
    END
  END w0_wd_in[279]
  PIN w0_wd_in[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 33.025 0.000 33.095 0.140 ;
    END
  END w0_wd_in[280]
  PIN w0_wd_in[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 34.355 0.000 34.425 0.140 ;
    END
  END w0_wd_in[281]
  PIN w0_wd_in[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 35.685 0.000 35.755 0.140 ;
    END
  END w0_wd_in[282]
  PIN w0_wd_in[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 37.015 0.000 37.085 0.140 ;
    END
  END w0_wd_in[283]
  PIN w0_wd_in[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 38.345 0.000 38.415 0.140 ;
    END
  END w0_wd_in[284]
  PIN w0_wd_in[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 39.675 0.000 39.745 0.140 ;
    END
  END w0_wd_in[285]
  PIN w0_wd_in[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 41.005 0.000 41.075 0.140 ;
    END
  END w0_wd_in[286]
  PIN w0_wd_in[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 42.335 0.000 42.405 0.140 ;
    END
  END w0_wd_in[287]
  PIN w0_wd_in[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 43.665 0.000 43.735 0.140 ;
    END
  END w0_wd_in[288]
  PIN w0_wd_in[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 44.995 0.000 45.065 0.140 ;
    END
  END w0_wd_in[289]
  PIN w0_wd_in[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 46.325 0.000 46.395 0.140 ;
    END
  END w0_wd_in[290]
  PIN w0_wd_in[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 47.655 0.000 47.725 0.140 ;
    END
  END w0_wd_in[291]
  PIN w0_wd_in[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 48.985 0.000 49.055 0.140 ;
    END
  END w0_wd_in[292]
  PIN w0_wd_in[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 50.315 0.000 50.385 0.140 ;
    END
  END w0_wd_in[293]
  PIN w0_wd_in[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 51.645 0.000 51.715 0.140 ;
    END
  END w0_wd_in[294]
  PIN w0_wd_in[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 52.975 0.000 53.045 0.140 ;
    END
  END w0_wd_in[295]
  PIN w0_wd_in[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 54.305 0.000 54.375 0.140 ;
    END
  END w0_wd_in[296]
  PIN w0_wd_in[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 55.635 0.000 55.705 0.140 ;
    END
  END w0_wd_in[297]
  PIN w0_wd_in[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 56.965 0.000 57.035 0.140 ;
    END
  END w0_wd_in[298]
  PIN w0_wd_in[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 58.295 0.000 58.365 0.140 ;
    END
  END w0_wd_in[299]
  PIN w0_wd_in[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 59.625 0.000 59.695 0.140 ;
    END
  END w0_wd_in[300]
  PIN w0_wd_in[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 60.955 0.000 61.025 0.140 ;
    END
  END w0_wd_in[301]
  PIN w0_wd_in[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 62.285 0.000 62.355 0.140 ;
    END
  END w0_wd_in[302]
  PIN w0_wd_in[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 63.615 0.000 63.685 0.140 ;
    END
  END w0_wd_in[303]
  PIN w0_wd_in[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 64.945 0.000 65.015 0.140 ;
    END
  END w0_wd_in[304]
  PIN w0_wd_in[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 66.275 0.000 66.345 0.140 ;
    END
  END w0_wd_in[305]
  PIN w0_wd_in[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 67.605 0.000 67.675 0.140 ;
    END
  END w0_wd_in[306]
  PIN w0_wd_in[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 68.935 0.000 69.005 0.140 ;
    END
  END w0_wd_in[307]
  PIN w0_wd_in[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 70.265 0.000 70.335 0.140 ;
    END
  END w0_wd_in[308]
  PIN w0_wd_in[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 71.595 0.000 71.665 0.140 ;
    END
  END w0_wd_in[309]
  PIN w0_wd_in[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 72.925 0.000 72.995 0.140 ;
    END
  END w0_wd_in[310]
  PIN w0_wd_in[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 74.255 0.000 74.325 0.140 ;
    END
  END w0_wd_in[311]
  PIN w0_wd_in[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 75.585 0.000 75.655 0.140 ;
    END
  END w0_wd_in[312]
  PIN w0_wd_in[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 76.915 0.000 76.985 0.140 ;
    END
  END w0_wd_in[313]
  PIN w0_wd_in[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 78.245 0.000 78.315 0.140 ;
    END
  END w0_wd_in[314]
  PIN w0_wd_in[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 79.575 0.000 79.645 0.140 ;
    END
  END w0_wd_in[315]
  PIN w0_wd_in[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 80.905 0.000 80.975 0.140 ;
    END
  END w0_wd_in[316]
  PIN w0_wd_in[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 82.235 0.000 82.305 0.140 ;
    END
  END w0_wd_in[317]
  PIN w0_wd_in[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 83.565 0.000 83.635 0.140 ;
    END
  END w0_wd_in[318]
  PIN w0_wd_in[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 84.895 0.000 84.965 0.140 ;
    END
  END w0_wd_in[319]
  PIN w0_wd_in[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 86.225 0.000 86.295 0.140 ;
    END
  END w0_wd_in[320]
  PIN w0_wd_in[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 87.555 0.000 87.625 0.140 ;
    END
  END w0_wd_in[321]
  PIN w0_wd_in[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 88.885 0.000 88.955 0.140 ;
    END
  END w0_wd_in[322]
  PIN w0_wd_in[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 90.215 0.000 90.285 0.140 ;
    END
  END w0_wd_in[323]
  PIN w0_wd_in[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 91.545 0.000 91.615 0.140 ;
    END
  END w0_wd_in[324]
  PIN w0_wd_in[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 92.875 0.000 92.945 0.140 ;
    END
  END w0_wd_in[325]
  PIN w0_wd_in[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 94.205 0.000 94.275 0.140 ;
    END
  END w0_wd_in[326]
  PIN w0_wd_in[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 95.535 0.000 95.605 0.140 ;
    END
  END w0_wd_in[327]
  PIN w0_wd_in[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 96.865 0.000 96.935 0.140 ;
    END
  END w0_wd_in[328]
  PIN w0_wd_in[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 98.195 0.000 98.265 0.140 ;
    END
  END w0_wd_in[329]
  PIN w0_wd_in[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 99.525 0.000 99.595 0.140 ;
    END
  END w0_wd_in[330]
  PIN w0_wd_in[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 100.855 0.000 100.925 0.140 ;
    END
  END w0_wd_in[331]
  PIN w0_wd_in[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 102.185 0.000 102.255 0.140 ;
    END
  END w0_wd_in[332]
  PIN w0_wd_in[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 103.515 0.000 103.585 0.140 ;
    END
  END w0_wd_in[333]
  PIN w0_wd_in[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 104.845 0.000 104.915 0.140 ;
    END
  END w0_wd_in[334]
  PIN w0_wd_in[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 106.175 0.000 106.245 0.140 ;
    END
  END w0_wd_in[335]
  PIN w0_wd_in[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 107.505 0.000 107.575 0.140 ;
    END
  END w0_wd_in[336]
  PIN w0_wd_in[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 108.835 0.000 108.905 0.140 ;
    END
  END w0_wd_in[337]
  PIN w0_wd_in[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 110.165 0.000 110.235 0.140 ;
    END
  END w0_wd_in[338]
  PIN w0_wd_in[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 111.495 0.000 111.565 0.140 ;
    END
  END w0_wd_in[339]
  PIN w0_wd_in[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 112.825 0.000 112.895 0.140 ;
    END
  END w0_wd_in[340]
  PIN w0_wd_in[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 114.155 0.000 114.225 0.140 ;
    END
  END w0_wd_in[341]
  PIN w0_wd_in[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 115.485 0.000 115.555 0.140 ;
    END
  END w0_wd_in[342]
  PIN w0_wd_in[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 116.815 0.000 116.885 0.140 ;
    END
  END w0_wd_in[343]
  PIN w0_wd_in[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 118.145 0.000 118.215 0.140 ;
    END
  END w0_wd_in[344]
  PIN w0_wd_in[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 119.475 0.000 119.545 0.140 ;
    END
  END w0_wd_in[345]
  PIN w0_wd_in[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 120.805 0.000 120.875 0.140 ;
    END
  END w0_wd_in[346]
  PIN w0_wd_in[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 122.135 0.000 122.205 0.140 ;
    END
  END w0_wd_in[347]
  PIN w0_wd_in[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 123.465 0.000 123.535 0.140 ;
    END
  END w0_wd_in[348]
  PIN w0_wd_in[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 124.795 0.000 124.865 0.140 ;
    END
  END w0_wd_in[349]
  PIN w0_wd_in[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 126.125 0.000 126.195 0.140 ;
    END
  END w0_wd_in[350]
  PIN w0_wd_in[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 127.455 0.000 127.525 0.140 ;
    END
  END w0_wd_in[351]
  PIN w0_wd_in[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 128.785 0.000 128.855 0.140 ;
    END
  END w0_wd_in[352]
  PIN w0_wd_in[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 130.115 0.000 130.185 0.140 ;
    END
  END w0_wd_in[353]
  PIN w0_wd_in[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 131.445 0.000 131.515 0.140 ;
    END
  END w0_wd_in[354]
  PIN w0_wd_in[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 132.775 0.000 132.845 0.140 ;
    END
  END w0_wd_in[355]
  PIN w0_wd_in[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 134.105 0.000 134.175 0.140 ;
    END
  END w0_wd_in[356]
  PIN w0_wd_in[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 135.435 0.000 135.505 0.140 ;
    END
  END w0_wd_in[357]
  PIN w0_wd_in[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 136.765 0.000 136.835 0.140 ;
    END
  END w0_wd_in[358]
  PIN w0_wd_in[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 138.095 0.000 138.165 0.140 ;
    END
  END w0_wd_in[359]
  PIN w0_wd_in[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 139.425 0.000 139.495 0.140 ;
    END
  END w0_wd_in[360]
  PIN w0_wd_in[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 140.755 0.000 140.825 0.140 ;
    END
  END w0_wd_in[361]
  PIN w0_wd_in[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 142.085 0.000 142.155 0.140 ;
    END
  END w0_wd_in[362]
  PIN w0_wd_in[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 143.415 0.000 143.485 0.140 ;
    END
  END w0_wd_in[363]
  PIN w0_wd_in[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 144.745 0.000 144.815 0.140 ;
    END
  END w0_wd_in[364]
  PIN w0_wd_in[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 146.075 0.000 146.145 0.140 ;
    END
  END w0_wd_in[365]
  PIN w0_wd_in[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 147.405 0.000 147.475 0.140 ;
    END
  END w0_wd_in[366]
  PIN w0_wd_in[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 148.735 0.000 148.805 0.140 ;
    END
  END w0_wd_in[367]
  PIN w0_wd_in[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 150.065 0.000 150.135 0.140 ;
    END
  END w0_wd_in[368]
  PIN w0_wd_in[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 151.395 0.000 151.465 0.140 ;
    END
  END w0_wd_in[369]
  PIN w0_wd_in[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 152.725 0.000 152.795 0.140 ;
    END
  END w0_wd_in[370]
  PIN w0_wd_in[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 154.055 0.000 154.125 0.140 ;
    END
  END w0_wd_in[371]
  PIN w0_wd_in[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 155.385 0.000 155.455 0.140 ;
    END
  END w0_wd_in[372]
  PIN w0_wd_in[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 156.715 0.000 156.785 0.140 ;
    END
  END w0_wd_in[373]
  PIN w0_wd_in[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 158.045 0.000 158.115 0.140 ;
    END
  END w0_wd_in[374]
  PIN w0_wd_in[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 159.375 0.000 159.445 0.140 ;
    END
  END w0_wd_in[375]
  PIN w0_wd_in[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 160.705 0.000 160.775 0.140 ;
    END
  END w0_wd_in[376]
  PIN w0_wd_in[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 162.035 0.000 162.105 0.140 ;
    END
  END w0_wd_in[377]
  PIN w0_wd_in[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 163.365 0.000 163.435 0.140 ;
    END
  END w0_wd_in[378]
  PIN w0_wd_in[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 164.695 0.000 164.765 0.140 ;
    END
  END w0_wd_in[379]
  PIN w0_wd_in[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 166.025 0.000 166.095 0.140 ;
    END
  END w0_wd_in[380]
  PIN w0_wd_in[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 167.355 0.000 167.425 0.140 ;
    END
  END w0_wd_in[381]
  PIN w0_wd_in[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 168.685 0.000 168.755 0.140 ;
    END
  END w0_wd_in[382]
  PIN w0_wd_in[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 170.015 0.000 170.085 0.140 ;
    END
  END w0_wd_in[383]
  PIN w0_wd_in[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 171.345 0.000 171.415 0.140 ;
    END
  END w0_wd_in[384]
  PIN w0_wd_in[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 172.675 0.000 172.745 0.140 ;
    END
  END w0_wd_in[385]
  PIN w0_wd_in[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 174.005 0.000 174.075 0.140 ;
    END
  END w0_wd_in[386]
  PIN w0_wd_in[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 175.335 0.000 175.405 0.140 ;
    END
  END w0_wd_in[387]
  PIN w0_wd_in[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 176.665 0.000 176.735 0.140 ;
    END
  END w0_wd_in[388]
  PIN w0_wd_in[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 177.995 0.000 178.065 0.140 ;
    END
  END w0_wd_in[389]
  PIN w0_wd_in[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 179.325 0.000 179.395 0.140 ;
    END
  END w0_wd_in[390]
  PIN w0_wd_in[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 180.655 0.000 180.725 0.140 ;
    END
  END w0_wd_in[391]
  PIN w0_wd_in[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 181.985 0.000 182.055 0.140 ;
    END
  END w0_wd_in[392]
  PIN w0_wd_in[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 183.315 0.000 183.385 0.140 ;
    END
  END w0_wd_in[393]
  PIN w0_wd_in[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 184.645 0.000 184.715 0.140 ;
    END
  END w0_wd_in[394]
  PIN w0_wd_in[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 185.975 0.000 186.045 0.140 ;
    END
  END w0_wd_in[395]
  PIN w0_wd_in[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 187.305 0.000 187.375 0.140 ;
    END
  END w0_wd_in[396]
  PIN w0_wd_in[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 188.635 0.000 188.705 0.140 ;
    END
  END w0_wd_in[397]
  PIN w0_wd_in[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 189.965 0.000 190.035 0.140 ;
    END
  END w0_wd_in[398]
  PIN w0_wd_in[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 191.295 0.000 191.365 0.140 ;
    END
  END w0_wd_in[399]
  PIN w0_wd_in[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 192.625 0.000 192.695 0.140 ;
    END
  END w0_wd_in[400]
  PIN w0_wd_in[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 193.955 0.000 194.025 0.140 ;
    END
  END w0_wd_in[401]
  PIN w0_wd_in[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 195.285 0.000 195.355 0.140 ;
    END
  END w0_wd_in[402]
  PIN w0_wd_in[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 196.615 0.000 196.685 0.140 ;
    END
  END w0_wd_in[403]
  PIN w0_wd_in[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 197.945 0.000 198.015 0.140 ;
    END
  END w0_wd_in[404]
  PIN w0_wd_in[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 199.275 0.000 199.345 0.140 ;
    END
  END w0_wd_in[405]
  PIN w0_wd_in[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 200.605 0.000 200.675 0.140 ;
    END
  END w0_wd_in[406]
  PIN w0_wd_in[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 201.935 0.000 202.005 0.140 ;
    END
  END w0_wd_in[407]
  PIN w0_wd_in[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 203.265 0.000 203.335 0.140 ;
    END
  END w0_wd_in[408]
  PIN w0_wd_in[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 204.595 0.000 204.665 0.140 ;
    END
  END w0_wd_in[409]
  PIN w0_wd_in[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 205.925 0.000 205.995 0.140 ;
    END
  END w0_wd_in[410]
  PIN w0_wd_in[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 207.255 0.000 207.325 0.140 ;
    END
  END w0_wd_in[411]
  PIN w0_wd_in[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 208.585 0.000 208.655 0.140 ;
    END
  END w0_wd_in[412]
  PIN w0_wd_in[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 209.915 0.000 209.985 0.140 ;
    END
  END w0_wd_in[413]
  PIN w0_wd_in[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 211.245 0.000 211.315 0.140 ;
    END
  END w0_wd_in[414]
  PIN w0_wd_in[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 212.575 0.000 212.645 0.140 ;
    END
  END w0_wd_in[415]
  PIN w0_wd_in[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 213.905 0.000 213.975 0.140 ;
    END
  END w0_wd_in[416]
  PIN w0_wd_in[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 215.235 0.000 215.305 0.140 ;
    END
  END w0_wd_in[417]
  PIN w0_wd_in[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 216.565 0.000 216.635 0.140 ;
    END
  END w0_wd_in[418]
  PIN w0_wd_in[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 217.895 0.000 217.965 0.140 ;
    END
  END w0_wd_in[419]
  PIN w0_wd_in[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 219.225 0.000 219.295 0.140 ;
    END
  END w0_wd_in[420]
  PIN w0_wd_in[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 220.555 0.000 220.625 0.140 ;
    END
  END w0_wd_in[421]
  PIN w0_wd_in[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 221.885 0.000 221.955 0.140 ;
    END
  END w0_wd_in[422]
  PIN w0_wd_in[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 223.215 0.000 223.285 0.140 ;
    END
  END w0_wd_in[423]
  PIN w0_wd_in[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 224.545 0.000 224.615 0.140 ;
    END
  END w0_wd_in[424]
  PIN w0_wd_in[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 225.875 0.000 225.945 0.140 ;
    END
  END w0_wd_in[425]
  PIN w0_wd_in[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 227.205 0.000 227.275 0.140 ;
    END
  END w0_wd_in[426]
  PIN w0_wd_in[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 228.535 0.000 228.605 0.140 ;
    END
  END w0_wd_in[427]
  PIN w0_wd_in[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 229.865 0.000 229.935 0.140 ;
    END
  END w0_wd_in[428]
  PIN w0_wd_in[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 231.195 0.000 231.265 0.140 ;
    END
  END w0_wd_in[429]
  PIN w0_wd_in[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 232.525 0.000 232.595 0.140 ;
    END
  END w0_wd_in[430]
  PIN w0_wd_in[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 233.855 0.000 233.925 0.140 ;
    END
  END w0_wd_in[431]
  PIN w0_wd_in[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 235.185 0.000 235.255 0.140 ;
    END
  END w0_wd_in[432]
  PIN w0_wd_in[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 236.515 0.000 236.585 0.140 ;
    END
  END w0_wd_in[433]
  PIN w0_wd_in[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 237.845 0.000 237.915 0.140 ;
    END
  END w0_wd_in[434]
  PIN w0_wd_in[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 239.175 0.000 239.245 0.140 ;
    END
  END w0_wd_in[435]
  PIN w0_wd_in[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 240.505 0.000 240.575 0.140 ;
    END
  END w0_wd_in[436]
  PIN w0_wd_in[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 241.835 0.000 241.905 0.140 ;
    END
  END w0_wd_in[437]
  PIN w0_wd_in[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 243.165 0.000 243.235 0.140 ;
    END
  END w0_wd_in[438]
  PIN w0_wd_in[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 244.495 0.000 244.565 0.140 ;
    END
  END w0_wd_in[439]
  PIN w0_wd_in[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 245.825 0.000 245.895 0.140 ;
    END
  END w0_wd_in[440]
  PIN w0_wd_in[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 247.155 0.000 247.225 0.140 ;
    END
  END w0_wd_in[441]
  PIN w0_wd_in[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 248.485 0.000 248.555 0.140 ;
    END
  END w0_wd_in[442]
  PIN w0_wd_in[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 249.815 0.000 249.885 0.140 ;
    END
  END w0_wd_in[443]
  PIN w0_wd_in[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 251.145 0.000 251.215 0.140 ;
    END
  END w0_wd_in[444]
  PIN w0_wd_in[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 252.475 0.000 252.545 0.140 ;
    END
  END w0_wd_in[445]
  PIN w0_wd_in[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 253.805 0.000 253.875 0.140 ;
    END
  END w0_wd_in[446]
  PIN w0_wd_in[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 255.135 0.000 255.205 0.140 ;
    END
  END w0_wd_in[447]
  PIN w0_wd_in[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 256.465 0.000 256.535 0.140 ;
    END
  END w0_wd_in[448]
  PIN w0_wd_in[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 257.795 0.000 257.865 0.140 ;
    END
  END w0_wd_in[449]
  PIN w0_wd_in[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 259.125 0.000 259.195 0.140 ;
    END
  END w0_wd_in[450]
  PIN w0_wd_in[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 260.455 0.000 260.525 0.140 ;
    END
  END w0_wd_in[451]
  PIN w0_wd_in[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 261.785 0.000 261.855 0.140 ;
    END
  END w0_wd_in[452]
  PIN w0_wd_in[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 263.115 0.000 263.185 0.140 ;
    END
  END w0_wd_in[453]
  PIN w0_wd_in[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 264.445 0.000 264.515 0.140 ;
    END
  END w0_wd_in[454]
  PIN w0_wd_in[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 265.775 0.000 265.845 0.140 ;
    END
  END w0_wd_in[455]
  PIN w0_wd_in[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 267.105 0.000 267.175 0.140 ;
    END
  END w0_wd_in[456]
  PIN w0_wd_in[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 268.435 0.000 268.505 0.140 ;
    END
  END w0_wd_in[457]
  PIN w0_wd_in[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 269.765 0.000 269.835 0.140 ;
    END
  END w0_wd_in[458]
  PIN w0_wd_in[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 271.095 0.000 271.165 0.140 ;
    END
  END w0_wd_in[459]
  PIN w0_wd_in[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 272.425 0.000 272.495 0.140 ;
    END
  END w0_wd_in[460]
  PIN w0_wd_in[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 273.755 0.000 273.825 0.140 ;
    END
  END w0_wd_in[461]
  PIN w0_wd_in[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 275.085 0.000 275.155 0.140 ;
    END
  END w0_wd_in[462]
  PIN w0_wd_in[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 276.415 0.000 276.485 0.140 ;
    END
  END w0_wd_in[463]
  PIN w0_wd_in[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 277.745 0.000 277.815 0.140 ;
    END
  END w0_wd_in[464]
  PIN w0_wd_in[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 279.075 0.000 279.145 0.140 ;
    END
  END w0_wd_in[465]
  PIN w0_wd_in[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 280.405 0.000 280.475 0.140 ;
    END
  END w0_wd_in[466]
  PIN w0_wd_in[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 281.735 0.000 281.805 0.140 ;
    END
  END w0_wd_in[467]
  PIN w0_wd_in[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 283.065 0.000 283.135 0.140 ;
    END
  END w0_wd_in[468]
  PIN w0_wd_in[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 284.395 0.000 284.465 0.140 ;
    END
  END w0_wd_in[469]
  PIN w0_wd_in[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 285.725 0.000 285.795 0.140 ;
    END
  END w0_wd_in[470]
  PIN w0_wd_in[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 287.055 0.000 287.125 0.140 ;
    END
  END w0_wd_in[471]
  PIN w0_wd_in[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 288.385 0.000 288.455 0.140 ;
    END
  END w0_wd_in[472]
  PIN w0_wd_in[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 289.715 0.000 289.785 0.140 ;
    END
  END w0_wd_in[473]
  PIN w0_wd_in[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 291.045 0.000 291.115 0.140 ;
    END
  END w0_wd_in[474]
  PIN w0_wd_in[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 292.375 0.000 292.445 0.140 ;
    END
  END w0_wd_in[475]
  PIN w0_wd_in[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 293.705 0.000 293.775 0.140 ;
    END
  END w0_wd_in[476]
  PIN w0_wd_in[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 295.035 0.000 295.105 0.140 ;
    END
  END w0_wd_in[477]
  PIN w0_wd_in[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 296.365 0.000 296.435 0.140 ;
    END
  END w0_wd_in[478]
  PIN w0_wd_in[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 297.695 0.000 297.765 0.140 ;
    END
  END w0_wd_in[479]
  PIN w0_wd_in[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 299.025 0.000 299.095 0.140 ;
    END
  END w0_wd_in[480]
  PIN w0_wd_in[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 300.355 0.000 300.425 0.140 ;
    END
  END w0_wd_in[481]
  PIN w0_wd_in[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 301.685 0.000 301.755 0.140 ;
    END
  END w0_wd_in[482]
  PIN w0_wd_in[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 303.015 0.000 303.085 0.140 ;
    END
  END w0_wd_in[483]
  PIN w0_wd_in[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 304.345 0.000 304.415 0.140 ;
    END
  END w0_wd_in[484]
  PIN w0_wd_in[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 305.675 0.000 305.745 0.140 ;
    END
  END w0_wd_in[485]
  PIN w0_wd_in[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 307.005 0.000 307.075 0.140 ;
    END
  END w0_wd_in[486]
  PIN w0_wd_in[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 308.335 0.000 308.405 0.140 ;
    END
  END w0_wd_in[487]
  PIN w0_wd_in[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 309.665 0.000 309.735 0.140 ;
    END
  END w0_wd_in[488]
  PIN w0_wd_in[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 310.995 0.000 311.065 0.140 ;
    END
  END w0_wd_in[489]
  PIN w0_wd_in[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 312.325 0.000 312.395 0.140 ;
    END
  END w0_wd_in[490]
  PIN w0_wd_in[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 313.655 0.000 313.725 0.140 ;
    END
  END w0_wd_in[491]
  PIN w0_wd_in[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 314.985 0.000 315.055 0.140 ;
    END
  END w0_wd_in[492]
  PIN w0_wd_in[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 316.315 0.000 316.385 0.140 ;
    END
  END w0_wd_in[493]
  PIN w0_wd_in[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 317.645 0.000 317.715 0.140 ;
    END
  END w0_wd_in[494]
  PIN w0_wd_in[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 318.975 0.000 319.045 0.140 ;
    END
  END w0_wd_in[495]
  PIN w0_wd_in[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 320.305 0.000 320.375 0.140 ;
    END
  END w0_wd_in[496]
  PIN w0_wd_in[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 321.635 0.000 321.705 0.140 ;
    END
  END w0_wd_in[497]
  PIN w0_wd_in[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 322.965 0.000 323.035 0.140 ;
    END
  END w0_wd_in[498]
  PIN w0_wd_in[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 324.295 0.000 324.365 0.140 ;
    END
  END w0_wd_in[499]
  PIN w0_wd_in[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 325.625 0.000 325.695 0.140 ;
    END
  END w0_wd_in[500]
  PIN w0_wd_in[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 326.955 0.000 327.025 0.140 ;
    END
  END w0_wd_in[501]
  PIN w0_wd_in[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 328.285 0.000 328.355 0.140 ;
    END
  END w0_wd_in[502]
  PIN w0_wd_in[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 329.615 0.000 329.685 0.140 ;
    END
  END w0_wd_in[503]
  PIN w0_wd_in[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 330.945 0.000 331.015 0.140 ;
    END
  END w0_wd_in[504]
  PIN w0_wd_in[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 332.275 0.000 332.345 0.140 ;
    END
  END w0_wd_in[505]
  PIN w0_wd_in[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 333.605 0.000 333.675 0.140 ;
    END
  END w0_wd_in[506]
  PIN w0_wd_in[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 334.935 0.000 335.005 0.140 ;
    END
  END w0_wd_in[507]
  PIN w0_wd_in[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 336.265 0.000 336.335 0.140 ;
    END
  END w0_wd_in[508]
  PIN w0_wd_in[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 337.595 0.000 337.665 0.140 ;
    END
  END w0_wd_in[509]
  PIN w0_wd_in[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 338.925 0.000 338.995 0.140 ;
    END
  END w0_wd_in[510]
  PIN w0_wd_in[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 340.255 0.000 340.325 0.140 ;
    END
  END w0_wd_in[511]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 341.585 0.000 341.655 0.140 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 342.915 0.000 342.985 0.140 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 344.245 0.000 344.315 0.140 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 345.575 0.000 345.645 0.140 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 346.905 0.000 346.975 0.140 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 348.235 0.000 348.305 0.140 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 349.565 0.000 349.635 0.140 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 350.895 0.000 350.965 0.140 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 352.225 0.000 352.295 0.140 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 353.555 0.000 353.625 0.140 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 354.885 0.000 354.955 0.140 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 356.215 0.000 356.285 0.140 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 357.545 0.000 357.615 0.140 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 358.875 0.000 358.945 0.140 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 360.205 0.000 360.275 0.140 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 361.535 0.000 361.605 0.140 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 362.865 0.000 362.935 0.140 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 364.195 0.000 364.265 0.140 ;
    END
  END r0_rd_out[17]
  PIN r0_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 365.525 0.000 365.595 0.140 ;
    END
  END r0_rd_out[18]
  PIN r0_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 366.855 0.000 366.925 0.140 ;
    END
  END r0_rd_out[19]
  PIN r0_rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 368.185 0.000 368.255 0.140 ;
    END
  END r0_rd_out[20]
  PIN r0_rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 369.515 0.000 369.585 0.140 ;
    END
  END r0_rd_out[21]
  PIN r0_rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 370.845 0.000 370.915 0.140 ;
    END
  END r0_rd_out[22]
  PIN r0_rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 372.175 0.000 372.245 0.140 ;
    END
  END r0_rd_out[23]
  PIN r0_rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 373.505 0.000 373.575 0.140 ;
    END
  END r0_rd_out[24]
  PIN r0_rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 374.835 0.000 374.905 0.140 ;
    END
  END r0_rd_out[25]
  PIN r0_rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 376.165 0.000 376.235 0.140 ;
    END
  END r0_rd_out[26]
  PIN r0_rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 377.495 0.000 377.565 0.140 ;
    END
  END r0_rd_out[27]
  PIN r0_rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 378.825 0.000 378.895 0.140 ;
    END
  END r0_rd_out[28]
  PIN r0_rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 380.155 0.000 380.225 0.140 ;
    END
  END r0_rd_out[29]
  PIN r0_rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 381.485 0.000 381.555 0.140 ;
    END
  END r0_rd_out[30]
  PIN r0_rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 382.815 0.000 382.885 0.140 ;
    END
  END r0_rd_out[31]
  PIN r0_rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 384.145 0.000 384.215 0.140 ;
    END
  END r0_rd_out[32]
  PIN r0_rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 385.475 0.000 385.545 0.140 ;
    END
  END r0_rd_out[33]
  PIN r0_rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 386.805 0.000 386.875 0.140 ;
    END
  END r0_rd_out[34]
  PIN r0_rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 388.135 0.000 388.205 0.140 ;
    END
  END r0_rd_out[35]
  PIN r0_rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 389.465 0.000 389.535 0.140 ;
    END
  END r0_rd_out[36]
  PIN r0_rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 390.795 0.000 390.865 0.140 ;
    END
  END r0_rd_out[37]
  PIN r0_rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 392.125 0.000 392.195 0.140 ;
    END
  END r0_rd_out[38]
  PIN r0_rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 393.455 0.000 393.525 0.140 ;
    END
  END r0_rd_out[39]
  PIN r0_rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 394.785 0.000 394.855 0.140 ;
    END
  END r0_rd_out[40]
  PIN r0_rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 396.115 0.000 396.185 0.140 ;
    END
  END r0_rd_out[41]
  PIN r0_rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 397.445 0.000 397.515 0.140 ;
    END
  END r0_rd_out[42]
  PIN r0_rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 398.775 0.000 398.845 0.140 ;
    END
  END r0_rd_out[43]
  PIN r0_rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 400.105 0.000 400.175 0.140 ;
    END
  END r0_rd_out[44]
  PIN r0_rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 401.435 0.000 401.505 0.140 ;
    END
  END r0_rd_out[45]
  PIN r0_rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 402.765 0.000 402.835 0.140 ;
    END
  END r0_rd_out[46]
  PIN r0_rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 404.095 0.000 404.165 0.140 ;
    END
  END r0_rd_out[47]
  PIN r0_rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 405.425 0.000 405.495 0.140 ;
    END
  END r0_rd_out[48]
  PIN r0_rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 406.755 0.000 406.825 0.140 ;
    END
  END r0_rd_out[49]
  PIN r0_rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 408.085 0.000 408.155 0.140 ;
    END
  END r0_rd_out[50]
  PIN r0_rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 409.415 0.000 409.485 0.140 ;
    END
  END r0_rd_out[51]
  PIN r0_rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 410.745 0.000 410.815 0.140 ;
    END
  END r0_rd_out[52]
  PIN r0_rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 412.075 0.000 412.145 0.140 ;
    END
  END r0_rd_out[53]
  PIN r0_rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 413.405 0.000 413.475 0.140 ;
    END
  END r0_rd_out[54]
  PIN r0_rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 414.735 0.000 414.805 0.140 ;
    END
  END r0_rd_out[55]
  PIN r0_rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 416.065 0.000 416.135 0.140 ;
    END
  END r0_rd_out[56]
  PIN r0_rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 417.395 0.000 417.465 0.140 ;
    END
  END r0_rd_out[57]
  PIN r0_rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 418.725 0.000 418.795 0.140 ;
    END
  END r0_rd_out[58]
  PIN r0_rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 420.055 0.000 420.125 0.140 ;
    END
  END r0_rd_out[59]
  PIN r0_rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 421.385 0.000 421.455 0.140 ;
    END
  END r0_rd_out[60]
  PIN r0_rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 422.715 0.000 422.785 0.140 ;
    END
  END r0_rd_out[61]
  PIN r0_rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 424.045 0.000 424.115 0.140 ;
    END
  END r0_rd_out[62]
  PIN r0_rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 425.375 0.000 425.445 0.140 ;
    END
  END r0_rd_out[63]
  PIN r0_rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 426.705 0.000 426.775 0.140 ;
    END
  END r0_rd_out[64]
  PIN r0_rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 428.035 0.000 428.105 0.140 ;
    END
  END r0_rd_out[65]
  PIN r0_rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 429.365 0.000 429.435 0.140 ;
    END
  END r0_rd_out[66]
  PIN r0_rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 430.695 0.000 430.765 0.140 ;
    END
  END r0_rd_out[67]
  PIN r0_rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 432.025 0.000 432.095 0.140 ;
    END
  END r0_rd_out[68]
  PIN r0_rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 433.355 0.000 433.425 0.140 ;
    END
  END r0_rd_out[69]
  PIN r0_rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 434.685 0.000 434.755 0.140 ;
    END
  END r0_rd_out[70]
  PIN r0_rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 436.015 0.000 436.085 0.140 ;
    END
  END r0_rd_out[71]
  PIN r0_rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 437.345 0.000 437.415 0.140 ;
    END
  END r0_rd_out[72]
  PIN r0_rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 438.675 0.000 438.745 0.140 ;
    END
  END r0_rd_out[73]
  PIN r0_rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 440.005 0.000 440.075 0.140 ;
    END
  END r0_rd_out[74]
  PIN r0_rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 441.335 0.000 441.405 0.140 ;
    END
  END r0_rd_out[75]
  PIN r0_rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 442.665 0.000 442.735 0.140 ;
    END
  END r0_rd_out[76]
  PIN r0_rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 443.995 0.000 444.065 0.140 ;
    END
  END r0_rd_out[77]
  PIN r0_rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 445.325 0.000 445.395 0.140 ;
    END
  END r0_rd_out[78]
  PIN r0_rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 446.655 0.000 446.725 0.140 ;
    END
  END r0_rd_out[79]
  PIN r0_rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 447.985 0.000 448.055 0.140 ;
    END
  END r0_rd_out[80]
  PIN r0_rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 449.315 0.000 449.385 0.140 ;
    END
  END r0_rd_out[81]
  PIN r0_rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 450.645 0.000 450.715 0.140 ;
    END
  END r0_rd_out[82]
  PIN r0_rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 451.975 0.000 452.045 0.140 ;
    END
  END r0_rd_out[83]
  PIN r0_rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 453.305 0.000 453.375 0.140 ;
    END
  END r0_rd_out[84]
  PIN r0_rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 454.635 0.000 454.705 0.140 ;
    END
  END r0_rd_out[85]
  PIN r0_rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 455.965 0.000 456.035 0.140 ;
    END
  END r0_rd_out[86]
  PIN r0_rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 457.295 0.000 457.365 0.140 ;
    END
  END r0_rd_out[87]
  PIN r0_rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 458.625 0.000 458.695 0.140 ;
    END
  END r0_rd_out[88]
  PIN r0_rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 459.955 0.000 460.025 0.140 ;
    END
  END r0_rd_out[89]
  PIN r0_rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 461.285 0.000 461.355 0.140 ;
    END
  END r0_rd_out[90]
  PIN r0_rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 462.615 0.000 462.685 0.140 ;
    END
  END r0_rd_out[91]
  PIN r0_rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 463.945 0.000 464.015 0.140 ;
    END
  END r0_rd_out[92]
  PIN r0_rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 465.275 0.000 465.345 0.140 ;
    END
  END r0_rd_out[93]
  PIN r0_rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 466.605 0.000 466.675 0.140 ;
    END
  END r0_rd_out[94]
  PIN r0_rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 467.935 0.000 468.005 0.140 ;
    END
  END r0_rd_out[95]
  PIN r0_rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 469.265 0.000 469.335 0.140 ;
    END
  END r0_rd_out[96]
  PIN r0_rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 470.595 0.000 470.665 0.140 ;
    END
  END r0_rd_out[97]
  PIN r0_rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 471.925 0.000 471.995 0.140 ;
    END
  END r0_rd_out[98]
  PIN r0_rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 473.255 0.000 473.325 0.140 ;
    END
  END r0_rd_out[99]
  PIN r0_rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 474.585 0.000 474.655 0.140 ;
    END
  END r0_rd_out[100]
  PIN r0_rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 475.915 0.000 475.985 0.140 ;
    END
  END r0_rd_out[101]
  PIN r0_rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 477.245 0.000 477.315 0.140 ;
    END
  END r0_rd_out[102]
  PIN r0_rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 478.575 0.000 478.645 0.140 ;
    END
  END r0_rd_out[103]
  PIN r0_rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 479.905 0.000 479.975 0.140 ;
    END
  END r0_rd_out[104]
  PIN r0_rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 481.235 0.000 481.305 0.140 ;
    END
  END r0_rd_out[105]
  PIN r0_rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 482.565 0.000 482.635 0.140 ;
    END
  END r0_rd_out[106]
  PIN r0_rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 483.895 0.000 483.965 0.140 ;
    END
  END r0_rd_out[107]
  PIN r0_rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 485.225 0.000 485.295 0.140 ;
    END
  END r0_rd_out[108]
  PIN r0_rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 486.555 0.000 486.625 0.140 ;
    END
  END r0_rd_out[109]
  PIN r0_rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 487.885 0.000 487.955 0.140 ;
    END
  END r0_rd_out[110]
  PIN r0_rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 489.215 0.000 489.285 0.140 ;
    END
  END r0_rd_out[111]
  PIN r0_rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 490.545 0.000 490.615 0.140 ;
    END
  END r0_rd_out[112]
  PIN r0_rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 491.875 0.000 491.945 0.140 ;
    END
  END r0_rd_out[113]
  PIN r0_rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 493.205 0.000 493.275 0.140 ;
    END
  END r0_rd_out[114]
  PIN r0_rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 494.535 0.000 494.605 0.140 ;
    END
  END r0_rd_out[115]
  PIN r0_rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 495.865 0.000 495.935 0.140 ;
    END
  END r0_rd_out[116]
  PIN r0_rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 497.195 0.000 497.265 0.140 ;
    END
  END r0_rd_out[117]
  PIN r0_rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 498.525 0.000 498.595 0.140 ;
    END
  END r0_rd_out[118]
  PIN r0_rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 499.855 0.000 499.925 0.140 ;
    END
  END r0_rd_out[119]
  PIN r0_rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 501.185 0.000 501.255 0.140 ;
    END
  END r0_rd_out[120]
  PIN r0_rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 502.515 0.000 502.585 0.140 ;
    END
  END r0_rd_out[121]
  PIN r0_rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 503.845 0.000 503.915 0.140 ;
    END
  END r0_rd_out[122]
  PIN r0_rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 505.175 0.000 505.245 0.140 ;
    END
  END r0_rd_out[123]
  PIN r0_rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 506.505 0.000 506.575 0.140 ;
    END
  END r0_rd_out[124]
  PIN r0_rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 507.835 0.000 507.905 0.140 ;
    END
  END r0_rd_out[125]
  PIN r0_rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 509.165 0.000 509.235 0.140 ;
    END
  END r0_rd_out[126]
  PIN r0_rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 510.495 0.000 510.565 0.140 ;
    END
  END r0_rd_out[127]
  PIN r0_rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 511.825 0.000 511.895 0.140 ;
    END
  END r0_rd_out[128]
  PIN r0_rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 513.155 0.000 513.225 0.140 ;
    END
  END r0_rd_out[129]
  PIN r0_rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 514.485 0.000 514.555 0.140 ;
    END
  END r0_rd_out[130]
  PIN r0_rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 515.815 0.000 515.885 0.140 ;
    END
  END r0_rd_out[131]
  PIN r0_rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 517.145 0.000 517.215 0.140 ;
    END
  END r0_rd_out[132]
  PIN r0_rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 518.475 0.000 518.545 0.140 ;
    END
  END r0_rd_out[133]
  PIN r0_rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 519.805 0.000 519.875 0.140 ;
    END
  END r0_rd_out[134]
  PIN r0_rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 521.135 0.000 521.205 0.140 ;
    END
  END r0_rd_out[135]
  PIN r0_rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 522.465 0.000 522.535 0.140 ;
    END
  END r0_rd_out[136]
  PIN r0_rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 523.795 0.000 523.865 0.140 ;
    END
  END r0_rd_out[137]
  PIN r0_rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 525.125 0.000 525.195 0.140 ;
    END
  END r0_rd_out[138]
  PIN r0_rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 526.455 0.000 526.525 0.140 ;
    END
  END r0_rd_out[139]
  PIN r0_rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 527.785 0.000 527.855 0.140 ;
    END
  END r0_rd_out[140]
  PIN r0_rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 529.115 0.000 529.185 0.140 ;
    END
  END r0_rd_out[141]
  PIN r0_rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 530.445 0.000 530.515 0.140 ;
    END
  END r0_rd_out[142]
  PIN r0_rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 531.775 0.000 531.845 0.140 ;
    END
  END r0_rd_out[143]
  PIN r0_rd_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 533.105 0.000 533.175 0.140 ;
    END
  END r0_rd_out[144]
  PIN r0_rd_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 534.435 0.000 534.505 0.140 ;
    END
  END r0_rd_out[145]
  PIN r0_rd_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 535.765 0.000 535.835 0.140 ;
    END
  END r0_rd_out[146]
  PIN r0_rd_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 537.095 0.000 537.165 0.140 ;
    END
  END r0_rd_out[147]
  PIN r0_rd_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 538.425 0.000 538.495 0.140 ;
    END
  END r0_rd_out[148]
  PIN r0_rd_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 539.755 0.000 539.825 0.140 ;
    END
  END r0_rd_out[149]
  PIN r0_rd_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 541.085 0.000 541.155 0.140 ;
    END
  END r0_rd_out[150]
  PIN r0_rd_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 542.415 0.000 542.485 0.140 ;
    END
  END r0_rd_out[151]
  PIN r0_rd_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 543.745 0.000 543.815 0.140 ;
    END
  END r0_rd_out[152]
  PIN r0_rd_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 545.075 0.000 545.145 0.140 ;
    END
  END r0_rd_out[153]
  PIN r0_rd_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 546.405 0.000 546.475 0.140 ;
    END
  END r0_rd_out[154]
  PIN r0_rd_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 547.735 0.000 547.805 0.140 ;
    END
  END r0_rd_out[155]
  PIN r0_rd_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 549.065 0.000 549.135 0.140 ;
    END
  END r0_rd_out[156]
  PIN r0_rd_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 550.395 0.000 550.465 0.140 ;
    END
  END r0_rd_out[157]
  PIN r0_rd_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 551.725 0.000 551.795 0.140 ;
    END
  END r0_rd_out[158]
  PIN r0_rd_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 553.055 0.000 553.125 0.140 ;
    END
  END r0_rd_out[159]
  PIN r0_rd_out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 554.385 0.000 554.455 0.140 ;
    END
  END r0_rd_out[160]
  PIN r0_rd_out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 555.715 0.000 555.785 0.140 ;
    END
  END r0_rd_out[161]
  PIN r0_rd_out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 557.045 0.000 557.115 0.140 ;
    END
  END r0_rd_out[162]
  PIN r0_rd_out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 558.375 0.000 558.445 0.140 ;
    END
  END r0_rd_out[163]
  PIN r0_rd_out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 559.705 0.000 559.775 0.140 ;
    END
  END r0_rd_out[164]
  PIN r0_rd_out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 561.035 0.000 561.105 0.140 ;
    END
  END r0_rd_out[165]
  PIN r0_rd_out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 562.365 0.000 562.435 0.140 ;
    END
  END r0_rd_out[166]
  PIN r0_rd_out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 563.695 0.000 563.765 0.140 ;
    END
  END r0_rd_out[167]
  PIN r0_rd_out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 565.025 0.000 565.095 0.140 ;
    END
  END r0_rd_out[168]
  PIN r0_rd_out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 566.355 0.000 566.425 0.140 ;
    END
  END r0_rd_out[169]
  PIN r0_rd_out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 567.685 0.000 567.755 0.140 ;
    END
  END r0_rd_out[170]
  PIN r0_rd_out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 569.015 0.000 569.085 0.140 ;
    END
  END r0_rd_out[171]
  PIN r0_rd_out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 570.345 0.000 570.415 0.140 ;
    END
  END r0_rd_out[172]
  PIN r0_rd_out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 571.675 0.000 571.745 0.140 ;
    END
  END r0_rd_out[173]
  PIN r0_rd_out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 573.005 0.000 573.075 0.140 ;
    END
  END r0_rd_out[174]
  PIN r0_rd_out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 574.335 0.000 574.405 0.140 ;
    END
  END r0_rd_out[175]
  PIN r0_rd_out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 575.665 0.000 575.735 0.140 ;
    END
  END r0_rd_out[176]
  PIN r0_rd_out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 576.995 0.000 577.065 0.140 ;
    END
  END r0_rd_out[177]
  PIN r0_rd_out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 578.325 0.000 578.395 0.140 ;
    END
  END r0_rd_out[178]
  PIN r0_rd_out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 579.655 0.000 579.725 0.140 ;
    END
  END r0_rd_out[179]
  PIN r0_rd_out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 580.985 0.000 581.055 0.140 ;
    END
  END r0_rd_out[180]
  PIN r0_rd_out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 582.315 0.000 582.385 0.140 ;
    END
  END r0_rd_out[181]
  PIN r0_rd_out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 583.645 0.000 583.715 0.140 ;
    END
  END r0_rd_out[182]
  PIN r0_rd_out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 584.975 0.000 585.045 0.140 ;
    END
  END r0_rd_out[183]
  PIN r0_rd_out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 586.305 0.000 586.375 0.140 ;
    END
  END r0_rd_out[184]
  PIN r0_rd_out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 587.635 0.000 587.705 0.140 ;
    END
  END r0_rd_out[185]
  PIN r0_rd_out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 588.965 0.000 589.035 0.140 ;
    END
  END r0_rd_out[186]
  PIN r0_rd_out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 590.295 0.000 590.365 0.140 ;
    END
  END r0_rd_out[187]
  PIN r0_rd_out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 591.625 0.000 591.695 0.140 ;
    END
  END r0_rd_out[188]
  PIN r0_rd_out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 592.955 0.000 593.025 0.140 ;
    END
  END r0_rd_out[189]
  PIN r0_rd_out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 594.285 0.000 594.355 0.140 ;
    END
  END r0_rd_out[190]
  PIN r0_rd_out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 595.615 0.000 595.685 0.140 ;
    END
  END r0_rd_out[191]
  PIN r0_rd_out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 596.945 0.000 597.015 0.140 ;
    END
  END r0_rd_out[192]
  PIN r0_rd_out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 598.275 0.000 598.345 0.140 ;
    END
  END r0_rd_out[193]
  PIN r0_rd_out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 599.605 0.000 599.675 0.140 ;
    END
  END r0_rd_out[194]
  PIN r0_rd_out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 600.935 0.000 601.005 0.140 ;
    END
  END r0_rd_out[195]
  PIN r0_rd_out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 602.265 0.000 602.335 0.140 ;
    END
  END r0_rd_out[196]
  PIN r0_rd_out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 603.595 0.000 603.665 0.140 ;
    END
  END r0_rd_out[197]
  PIN r0_rd_out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 604.925 0.000 604.995 0.140 ;
    END
  END r0_rd_out[198]
  PIN r0_rd_out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 606.255 0.000 606.325 0.140 ;
    END
  END r0_rd_out[199]
  PIN r0_rd_out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 607.585 0.000 607.655 0.140 ;
    END
  END r0_rd_out[200]
  PIN r0_rd_out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 608.915 0.000 608.985 0.140 ;
    END
  END r0_rd_out[201]
  PIN r0_rd_out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 610.245 0.000 610.315 0.140 ;
    END
  END r0_rd_out[202]
  PIN r0_rd_out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 611.575 0.000 611.645 0.140 ;
    END
  END r0_rd_out[203]
  PIN r0_rd_out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 612.905 0.000 612.975 0.140 ;
    END
  END r0_rd_out[204]
  PIN r0_rd_out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 614.235 0.000 614.305 0.140 ;
    END
  END r0_rd_out[205]
  PIN r0_rd_out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 615.565 0.000 615.635 0.140 ;
    END
  END r0_rd_out[206]
  PIN r0_rd_out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 616.895 0.000 616.965 0.140 ;
    END
  END r0_rd_out[207]
  PIN r0_rd_out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 618.225 0.000 618.295 0.140 ;
    END
  END r0_rd_out[208]
  PIN r0_rd_out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 619.555 0.000 619.625 0.140 ;
    END
  END r0_rd_out[209]
  PIN r0_rd_out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 620.885 0.000 620.955 0.140 ;
    END
  END r0_rd_out[210]
  PIN r0_rd_out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 622.215 0.000 622.285 0.140 ;
    END
  END r0_rd_out[211]
  PIN r0_rd_out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 623.545 0.000 623.615 0.140 ;
    END
  END r0_rd_out[212]
  PIN r0_rd_out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 624.875 0.000 624.945 0.140 ;
    END
  END r0_rd_out[213]
  PIN r0_rd_out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 626.205 0.000 626.275 0.140 ;
    END
  END r0_rd_out[214]
  PIN r0_rd_out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 627.535 0.000 627.605 0.140 ;
    END
  END r0_rd_out[215]
  PIN r0_rd_out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 628.865 0.000 628.935 0.140 ;
    END
  END r0_rd_out[216]
  PIN r0_rd_out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 630.195 0.000 630.265 0.140 ;
    END
  END r0_rd_out[217]
  PIN r0_rd_out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 631.525 0.000 631.595 0.140 ;
    END
  END r0_rd_out[218]
  PIN r0_rd_out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 632.855 0.000 632.925 0.140 ;
    END
  END r0_rd_out[219]
  PIN r0_rd_out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 634.185 0.000 634.255 0.140 ;
    END
  END r0_rd_out[220]
  PIN r0_rd_out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 635.515 0.000 635.585 0.140 ;
    END
  END r0_rd_out[221]
  PIN r0_rd_out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 636.845 0.000 636.915 0.140 ;
    END
  END r0_rd_out[222]
  PIN r0_rd_out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 638.175 0.000 638.245 0.140 ;
    END
  END r0_rd_out[223]
  PIN r0_rd_out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 639.505 0.000 639.575 0.140 ;
    END
  END r0_rd_out[224]
  PIN r0_rd_out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 640.835 0.000 640.905 0.140 ;
    END
  END r0_rd_out[225]
  PIN r0_rd_out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 642.165 0.000 642.235 0.140 ;
    END
  END r0_rd_out[226]
  PIN r0_rd_out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 643.495 0.000 643.565 0.140 ;
    END
  END r0_rd_out[227]
  PIN r0_rd_out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 644.825 0.000 644.895 0.140 ;
    END
  END r0_rd_out[228]
  PIN r0_rd_out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 646.155 0.000 646.225 0.140 ;
    END
  END r0_rd_out[229]
  PIN r0_rd_out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 647.485 0.000 647.555 0.140 ;
    END
  END r0_rd_out[230]
  PIN r0_rd_out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 648.815 0.000 648.885 0.140 ;
    END
  END r0_rd_out[231]
  PIN r0_rd_out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 650.145 0.000 650.215 0.140 ;
    END
  END r0_rd_out[232]
  PIN r0_rd_out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 651.475 0.000 651.545 0.140 ;
    END
  END r0_rd_out[233]
  PIN r0_rd_out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 652.805 0.000 652.875 0.140 ;
    END
  END r0_rd_out[234]
  PIN r0_rd_out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 654.135 0.000 654.205 0.140 ;
    END
  END r0_rd_out[235]
  PIN r0_rd_out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 655.465 0.000 655.535 0.140 ;
    END
  END r0_rd_out[236]
  PIN r0_rd_out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 656.795 0.000 656.865 0.140 ;
    END
  END r0_rd_out[237]
  PIN r0_rd_out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 658.125 0.000 658.195 0.140 ;
    END
  END r0_rd_out[238]
  PIN r0_rd_out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 659.455 0.000 659.525 0.140 ;
    END
  END r0_rd_out[239]
  PIN r0_rd_out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 660.785 0.000 660.855 0.140 ;
    END
  END r0_rd_out[240]
  PIN r0_rd_out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 662.115 0.000 662.185 0.140 ;
    END
  END r0_rd_out[241]
  PIN r0_rd_out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 663.445 0.000 663.515 0.140 ;
    END
  END r0_rd_out[242]
  PIN r0_rd_out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 664.775 0.000 664.845 0.140 ;
    END
  END r0_rd_out[243]
  PIN r0_rd_out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 666.105 0.000 666.175 0.140 ;
    END
  END r0_rd_out[244]
  PIN r0_rd_out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 667.435 0.000 667.505 0.140 ;
    END
  END r0_rd_out[245]
  PIN r0_rd_out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 668.765 0.000 668.835 0.140 ;
    END
  END r0_rd_out[246]
  PIN r0_rd_out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 670.095 0.000 670.165 0.140 ;
    END
  END r0_rd_out[247]
  PIN r0_rd_out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 671.425 0.000 671.495 0.140 ;
    END
  END r0_rd_out[248]
  PIN r0_rd_out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 672.755 0.000 672.825 0.140 ;
    END
  END r0_rd_out[249]
  PIN r0_rd_out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 674.085 0.000 674.155 0.140 ;
    END
  END r0_rd_out[250]
  PIN r0_rd_out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 675.415 0.000 675.485 0.140 ;
    END
  END r0_rd_out[251]
  PIN r0_rd_out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 676.745 0.000 676.815 0.140 ;
    END
  END r0_rd_out[252]
  PIN r0_rd_out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 678.075 0.000 678.145 0.140 ;
    END
  END r0_rd_out[253]
  PIN r0_rd_out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 679.405 0.000 679.475 0.140 ;
    END
  END r0_rd_out[254]
  PIN r0_rd_out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 680.735 0.000 680.805 0.140 ;
    END
  END r0_rd_out[255]
  PIN r0_rd_out[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1.105 767.060 1.175 767.200 ;
    END
  END r0_rd_out[256]
  PIN r0_rd_out[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 3.575 767.060 3.645 767.200 ;
    END
  END r0_rd_out[257]
  PIN r0_rd_out[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 6.045 767.060 6.115 767.200 ;
    END
  END r0_rd_out[258]
  PIN r0_rd_out[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 8.515 767.060 8.585 767.200 ;
    END
  END r0_rd_out[259]
  PIN r0_rd_out[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 10.985 767.060 11.055 767.200 ;
    END
  END r0_rd_out[260]
  PIN r0_rd_out[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 13.455 767.060 13.525 767.200 ;
    END
  END r0_rd_out[261]
  PIN r0_rd_out[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 15.925 767.060 15.995 767.200 ;
    END
  END r0_rd_out[262]
  PIN r0_rd_out[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 18.395 767.060 18.465 767.200 ;
    END
  END r0_rd_out[263]
  PIN r0_rd_out[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 20.865 767.060 20.935 767.200 ;
    END
  END r0_rd_out[264]
  PIN r0_rd_out[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 23.335 767.060 23.405 767.200 ;
    END
  END r0_rd_out[265]
  PIN r0_rd_out[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 25.805 767.060 25.875 767.200 ;
    END
  END r0_rd_out[266]
  PIN r0_rd_out[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 28.275 767.060 28.345 767.200 ;
    END
  END r0_rd_out[267]
  PIN r0_rd_out[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 30.745 767.060 30.815 767.200 ;
    END
  END r0_rd_out[268]
  PIN r0_rd_out[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 33.215 767.060 33.285 767.200 ;
    END
  END r0_rd_out[269]
  PIN r0_rd_out[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 35.685 767.060 35.755 767.200 ;
    END
  END r0_rd_out[270]
  PIN r0_rd_out[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 38.155 767.060 38.225 767.200 ;
    END
  END r0_rd_out[271]
  PIN r0_rd_out[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 40.625 767.060 40.695 767.200 ;
    END
  END r0_rd_out[272]
  PIN r0_rd_out[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 43.095 767.060 43.165 767.200 ;
    END
  END r0_rd_out[273]
  PIN r0_rd_out[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 45.565 767.060 45.635 767.200 ;
    END
  END r0_rd_out[274]
  PIN r0_rd_out[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 48.035 767.060 48.105 767.200 ;
    END
  END r0_rd_out[275]
  PIN r0_rd_out[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 50.505 767.060 50.575 767.200 ;
    END
  END r0_rd_out[276]
  PIN r0_rd_out[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 52.975 767.060 53.045 767.200 ;
    END
  END r0_rd_out[277]
  PIN r0_rd_out[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 55.445 767.060 55.515 767.200 ;
    END
  END r0_rd_out[278]
  PIN r0_rd_out[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 57.915 767.060 57.985 767.200 ;
    END
  END r0_rd_out[279]
  PIN r0_rd_out[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 60.385 767.060 60.455 767.200 ;
    END
  END r0_rd_out[280]
  PIN r0_rd_out[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 62.855 767.060 62.925 767.200 ;
    END
  END r0_rd_out[281]
  PIN r0_rd_out[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 65.325 767.060 65.395 767.200 ;
    END
  END r0_rd_out[282]
  PIN r0_rd_out[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 67.795 767.060 67.865 767.200 ;
    END
  END r0_rd_out[283]
  PIN r0_rd_out[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 70.265 767.060 70.335 767.200 ;
    END
  END r0_rd_out[284]
  PIN r0_rd_out[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 72.735 767.060 72.805 767.200 ;
    END
  END r0_rd_out[285]
  PIN r0_rd_out[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 75.205 767.060 75.275 767.200 ;
    END
  END r0_rd_out[286]
  PIN r0_rd_out[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 77.675 767.060 77.745 767.200 ;
    END
  END r0_rd_out[287]
  PIN r0_rd_out[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 80.145 767.060 80.215 767.200 ;
    END
  END r0_rd_out[288]
  PIN r0_rd_out[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 82.615 767.060 82.685 767.200 ;
    END
  END r0_rd_out[289]
  PIN r0_rd_out[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 85.085 767.060 85.155 767.200 ;
    END
  END r0_rd_out[290]
  PIN r0_rd_out[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 87.555 767.060 87.625 767.200 ;
    END
  END r0_rd_out[291]
  PIN r0_rd_out[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 90.025 767.060 90.095 767.200 ;
    END
  END r0_rd_out[292]
  PIN r0_rd_out[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 92.495 767.060 92.565 767.200 ;
    END
  END r0_rd_out[293]
  PIN r0_rd_out[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 94.965 767.060 95.035 767.200 ;
    END
  END r0_rd_out[294]
  PIN r0_rd_out[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 97.435 767.060 97.505 767.200 ;
    END
  END r0_rd_out[295]
  PIN r0_rd_out[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 99.905 767.060 99.975 767.200 ;
    END
  END r0_rd_out[296]
  PIN r0_rd_out[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 102.375 767.060 102.445 767.200 ;
    END
  END r0_rd_out[297]
  PIN r0_rd_out[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 104.845 767.060 104.915 767.200 ;
    END
  END r0_rd_out[298]
  PIN r0_rd_out[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 107.315 767.060 107.385 767.200 ;
    END
  END r0_rd_out[299]
  PIN r0_rd_out[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 109.785 767.060 109.855 767.200 ;
    END
  END r0_rd_out[300]
  PIN r0_rd_out[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 112.255 767.060 112.325 767.200 ;
    END
  END r0_rd_out[301]
  PIN r0_rd_out[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 114.725 767.060 114.795 767.200 ;
    END
  END r0_rd_out[302]
  PIN r0_rd_out[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 117.195 767.060 117.265 767.200 ;
    END
  END r0_rd_out[303]
  PIN r0_rd_out[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 119.665 767.060 119.735 767.200 ;
    END
  END r0_rd_out[304]
  PIN r0_rd_out[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 122.135 767.060 122.205 767.200 ;
    END
  END r0_rd_out[305]
  PIN r0_rd_out[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 124.605 767.060 124.675 767.200 ;
    END
  END r0_rd_out[306]
  PIN r0_rd_out[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 127.075 767.060 127.145 767.200 ;
    END
  END r0_rd_out[307]
  PIN r0_rd_out[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 129.545 767.060 129.615 767.200 ;
    END
  END r0_rd_out[308]
  PIN r0_rd_out[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 132.015 767.060 132.085 767.200 ;
    END
  END r0_rd_out[309]
  PIN r0_rd_out[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 134.485 767.060 134.555 767.200 ;
    END
  END r0_rd_out[310]
  PIN r0_rd_out[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 136.955 767.060 137.025 767.200 ;
    END
  END r0_rd_out[311]
  PIN r0_rd_out[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 139.425 767.060 139.495 767.200 ;
    END
  END r0_rd_out[312]
  PIN r0_rd_out[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 141.895 767.060 141.965 767.200 ;
    END
  END r0_rd_out[313]
  PIN r0_rd_out[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 144.365 767.060 144.435 767.200 ;
    END
  END r0_rd_out[314]
  PIN r0_rd_out[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 146.835 767.060 146.905 767.200 ;
    END
  END r0_rd_out[315]
  PIN r0_rd_out[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 149.305 767.060 149.375 767.200 ;
    END
  END r0_rd_out[316]
  PIN r0_rd_out[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 151.775 767.060 151.845 767.200 ;
    END
  END r0_rd_out[317]
  PIN r0_rd_out[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 154.245 767.060 154.315 767.200 ;
    END
  END r0_rd_out[318]
  PIN r0_rd_out[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 156.715 767.060 156.785 767.200 ;
    END
  END r0_rd_out[319]
  PIN r0_rd_out[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 159.185 767.060 159.255 767.200 ;
    END
  END r0_rd_out[320]
  PIN r0_rd_out[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 161.655 767.060 161.725 767.200 ;
    END
  END r0_rd_out[321]
  PIN r0_rd_out[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 164.125 767.060 164.195 767.200 ;
    END
  END r0_rd_out[322]
  PIN r0_rd_out[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 166.595 767.060 166.665 767.200 ;
    END
  END r0_rd_out[323]
  PIN r0_rd_out[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 169.065 767.060 169.135 767.200 ;
    END
  END r0_rd_out[324]
  PIN r0_rd_out[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 171.535 767.060 171.605 767.200 ;
    END
  END r0_rd_out[325]
  PIN r0_rd_out[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 174.005 767.060 174.075 767.200 ;
    END
  END r0_rd_out[326]
  PIN r0_rd_out[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 176.475 767.060 176.545 767.200 ;
    END
  END r0_rd_out[327]
  PIN r0_rd_out[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 178.945 767.060 179.015 767.200 ;
    END
  END r0_rd_out[328]
  PIN r0_rd_out[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 181.415 767.060 181.485 767.200 ;
    END
  END r0_rd_out[329]
  PIN r0_rd_out[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 183.885 767.060 183.955 767.200 ;
    END
  END r0_rd_out[330]
  PIN r0_rd_out[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 186.355 767.060 186.425 767.200 ;
    END
  END r0_rd_out[331]
  PIN r0_rd_out[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 188.825 767.060 188.895 767.200 ;
    END
  END r0_rd_out[332]
  PIN r0_rd_out[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 191.295 767.060 191.365 767.200 ;
    END
  END r0_rd_out[333]
  PIN r0_rd_out[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 193.765 767.060 193.835 767.200 ;
    END
  END r0_rd_out[334]
  PIN r0_rd_out[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 196.235 767.060 196.305 767.200 ;
    END
  END r0_rd_out[335]
  PIN r0_rd_out[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 198.705 767.060 198.775 767.200 ;
    END
  END r0_rd_out[336]
  PIN r0_rd_out[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 201.175 767.060 201.245 767.200 ;
    END
  END r0_rd_out[337]
  PIN r0_rd_out[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 203.645 767.060 203.715 767.200 ;
    END
  END r0_rd_out[338]
  PIN r0_rd_out[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 206.115 767.060 206.185 767.200 ;
    END
  END r0_rd_out[339]
  PIN r0_rd_out[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 208.585 767.060 208.655 767.200 ;
    END
  END r0_rd_out[340]
  PIN r0_rd_out[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 211.055 767.060 211.125 767.200 ;
    END
  END r0_rd_out[341]
  PIN r0_rd_out[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 213.525 767.060 213.595 767.200 ;
    END
  END r0_rd_out[342]
  PIN r0_rd_out[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 215.995 767.060 216.065 767.200 ;
    END
  END r0_rd_out[343]
  PIN r0_rd_out[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 218.465 767.060 218.535 767.200 ;
    END
  END r0_rd_out[344]
  PIN r0_rd_out[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 220.935 767.060 221.005 767.200 ;
    END
  END r0_rd_out[345]
  PIN r0_rd_out[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 223.405 767.060 223.475 767.200 ;
    END
  END r0_rd_out[346]
  PIN r0_rd_out[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 225.875 767.060 225.945 767.200 ;
    END
  END r0_rd_out[347]
  PIN r0_rd_out[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 228.345 767.060 228.415 767.200 ;
    END
  END r0_rd_out[348]
  PIN r0_rd_out[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 230.815 767.060 230.885 767.200 ;
    END
  END r0_rd_out[349]
  PIN r0_rd_out[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 233.285 767.060 233.355 767.200 ;
    END
  END r0_rd_out[350]
  PIN r0_rd_out[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 235.755 767.060 235.825 767.200 ;
    END
  END r0_rd_out[351]
  PIN r0_rd_out[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 238.225 767.060 238.295 767.200 ;
    END
  END r0_rd_out[352]
  PIN r0_rd_out[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 240.695 767.060 240.765 767.200 ;
    END
  END r0_rd_out[353]
  PIN r0_rd_out[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 243.165 767.060 243.235 767.200 ;
    END
  END r0_rd_out[354]
  PIN r0_rd_out[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 245.635 767.060 245.705 767.200 ;
    END
  END r0_rd_out[355]
  PIN r0_rd_out[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 248.105 767.060 248.175 767.200 ;
    END
  END r0_rd_out[356]
  PIN r0_rd_out[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 250.575 767.060 250.645 767.200 ;
    END
  END r0_rd_out[357]
  PIN r0_rd_out[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 253.045 767.060 253.115 767.200 ;
    END
  END r0_rd_out[358]
  PIN r0_rd_out[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 255.515 767.060 255.585 767.200 ;
    END
  END r0_rd_out[359]
  PIN r0_rd_out[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 257.985 767.060 258.055 767.200 ;
    END
  END r0_rd_out[360]
  PIN r0_rd_out[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 260.455 767.060 260.525 767.200 ;
    END
  END r0_rd_out[361]
  PIN r0_rd_out[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 262.925 767.060 262.995 767.200 ;
    END
  END r0_rd_out[362]
  PIN r0_rd_out[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 265.395 767.060 265.465 767.200 ;
    END
  END r0_rd_out[363]
  PIN r0_rd_out[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 267.865 767.060 267.935 767.200 ;
    END
  END r0_rd_out[364]
  PIN r0_rd_out[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 270.335 767.060 270.405 767.200 ;
    END
  END r0_rd_out[365]
  PIN r0_rd_out[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 272.805 767.060 272.875 767.200 ;
    END
  END r0_rd_out[366]
  PIN r0_rd_out[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 275.275 767.060 275.345 767.200 ;
    END
  END r0_rd_out[367]
  PIN r0_rd_out[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 277.745 767.060 277.815 767.200 ;
    END
  END r0_rd_out[368]
  PIN r0_rd_out[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 280.215 767.060 280.285 767.200 ;
    END
  END r0_rd_out[369]
  PIN r0_rd_out[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 282.685 767.060 282.755 767.200 ;
    END
  END r0_rd_out[370]
  PIN r0_rd_out[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 285.155 767.060 285.225 767.200 ;
    END
  END r0_rd_out[371]
  PIN r0_rd_out[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 287.625 767.060 287.695 767.200 ;
    END
  END r0_rd_out[372]
  PIN r0_rd_out[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 290.095 767.060 290.165 767.200 ;
    END
  END r0_rd_out[373]
  PIN r0_rd_out[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 292.565 767.060 292.635 767.200 ;
    END
  END r0_rd_out[374]
  PIN r0_rd_out[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 295.035 767.060 295.105 767.200 ;
    END
  END r0_rd_out[375]
  PIN r0_rd_out[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 297.505 767.060 297.575 767.200 ;
    END
  END r0_rd_out[376]
  PIN r0_rd_out[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 299.975 767.060 300.045 767.200 ;
    END
  END r0_rd_out[377]
  PIN r0_rd_out[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 302.445 767.060 302.515 767.200 ;
    END
  END r0_rd_out[378]
  PIN r0_rd_out[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 304.915 767.060 304.985 767.200 ;
    END
  END r0_rd_out[379]
  PIN r0_rd_out[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 307.385 767.060 307.455 767.200 ;
    END
  END r0_rd_out[380]
  PIN r0_rd_out[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 309.855 767.060 309.925 767.200 ;
    END
  END r0_rd_out[381]
  PIN r0_rd_out[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 312.325 767.060 312.395 767.200 ;
    END
  END r0_rd_out[382]
  PIN r0_rd_out[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 314.795 767.060 314.865 767.200 ;
    END
  END r0_rd_out[383]
  PIN r0_rd_out[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 317.265 767.060 317.335 767.200 ;
    END
  END r0_rd_out[384]
  PIN r0_rd_out[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 319.735 767.060 319.805 767.200 ;
    END
  END r0_rd_out[385]
  PIN r0_rd_out[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 322.205 767.060 322.275 767.200 ;
    END
  END r0_rd_out[386]
  PIN r0_rd_out[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 324.675 767.060 324.745 767.200 ;
    END
  END r0_rd_out[387]
  PIN r0_rd_out[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 327.145 767.060 327.215 767.200 ;
    END
  END r0_rd_out[388]
  PIN r0_rd_out[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 329.615 767.060 329.685 767.200 ;
    END
  END r0_rd_out[389]
  PIN r0_rd_out[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 332.085 767.060 332.155 767.200 ;
    END
  END r0_rd_out[390]
  PIN r0_rd_out[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 334.555 767.060 334.625 767.200 ;
    END
  END r0_rd_out[391]
  PIN r0_rd_out[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 337.025 767.060 337.095 767.200 ;
    END
  END r0_rd_out[392]
  PIN r0_rd_out[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 339.495 767.060 339.565 767.200 ;
    END
  END r0_rd_out[393]
  PIN r0_rd_out[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 341.965 767.060 342.035 767.200 ;
    END
  END r0_rd_out[394]
  PIN r0_rd_out[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 344.435 767.060 344.505 767.200 ;
    END
  END r0_rd_out[395]
  PIN r0_rd_out[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 346.905 767.060 346.975 767.200 ;
    END
  END r0_rd_out[396]
  PIN r0_rd_out[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 349.375 767.060 349.445 767.200 ;
    END
  END r0_rd_out[397]
  PIN r0_rd_out[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 351.845 767.060 351.915 767.200 ;
    END
  END r0_rd_out[398]
  PIN r0_rd_out[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 354.315 767.060 354.385 767.200 ;
    END
  END r0_rd_out[399]
  PIN r0_rd_out[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 356.785 767.060 356.855 767.200 ;
    END
  END r0_rd_out[400]
  PIN r0_rd_out[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 359.255 767.060 359.325 767.200 ;
    END
  END r0_rd_out[401]
  PIN r0_rd_out[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 361.725 767.060 361.795 767.200 ;
    END
  END r0_rd_out[402]
  PIN r0_rd_out[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 364.195 767.060 364.265 767.200 ;
    END
  END r0_rd_out[403]
  PIN r0_rd_out[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 366.665 767.060 366.735 767.200 ;
    END
  END r0_rd_out[404]
  PIN r0_rd_out[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 369.135 767.060 369.205 767.200 ;
    END
  END r0_rd_out[405]
  PIN r0_rd_out[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 371.605 767.060 371.675 767.200 ;
    END
  END r0_rd_out[406]
  PIN r0_rd_out[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 374.075 767.060 374.145 767.200 ;
    END
  END r0_rd_out[407]
  PIN r0_rd_out[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 376.545 767.060 376.615 767.200 ;
    END
  END r0_rd_out[408]
  PIN r0_rd_out[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 379.015 767.060 379.085 767.200 ;
    END
  END r0_rd_out[409]
  PIN r0_rd_out[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 381.485 767.060 381.555 767.200 ;
    END
  END r0_rd_out[410]
  PIN r0_rd_out[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 383.955 767.060 384.025 767.200 ;
    END
  END r0_rd_out[411]
  PIN r0_rd_out[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 386.425 767.060 386.495 767.200 ;
    END
  END r0_rd_out[412]
  PIN r0_rd_out[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 388.895 767.060 388.965 767.200 ;
    END
  END r0_rd_out[413]
  PIN r0_rd_out[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 391.365 767.060 391.435 767.200 ;
    END
  END r0_rd_out[414]
  PIN r0_rd_out[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 393.835 767.060 393.905 767.200 ;
    END
  END r0_rd_out[415]
  PIN r0_rd_out[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 396.305 767.060 396.375 767.200 ;
    END
  END r0_rd_out[416]
  PIN r0_rd_out[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 398.775 767.060 398.845 767.200 ;
    END
  END r0_rd_out[417]
  PIN r0_rd_out[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 401.245 767.060 401.315 767.200 ;
    END
  END r0_rd_out[418]
  PIN r0_rd_out[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 403.715 767.060 403.785 767.200 ;
    END
  END r0_rd_out[419]
  PIN r0_rd_out[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 406.185 767.060 406.255 767.200 ;
    END
  END r0_rd_out[420]
  PIN r0_rd_out[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 408.655 767.060 408.725 767.200 ;
    END
  END r0_rd_out[421]
  PIN r0_rd_out[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 411.125 767.060 411.195 767.200 ;
    END
  END r0_rd_out[422]
  PIN r0_rd_out[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 413.595 767.060 413.665 767.200 ;
    END
  END r0_rd_out[423]
  PIN r0_rd_out[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 416.065 767.060 416.135 767.200 ;
    END
  END r0_rd_out[424]
  PIN r0_rd_out[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 418.535 767.060 418.605 767.200 ;
    END
  END r0_rd_out[425]
  PIN r0_rd_out[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 421.005 767.060 421.075 767.200 ;
    END
  END r0_rd_out[426]
  PIN r0_rd_out[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 423.475 767.060 423.545 767.200 ;
    END
  END r0_rd_out[427]
  PIN r0_rd_out[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 425.945 767.060 426.015 767.200 ;
    END
  END r0_rd_out[428]
  PIN r0_rd_out[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 428.415 767.060 428.485 767.200 ;
    END
  END r0_rd_out[429]
  PIN r0_rd_out[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 430.885 767.060 430.955 767.200 ;
    END
  END r0_rd_out[430]
  PIN r0_rd_out[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 433.355 767.060 433.425 767.200 ;
    END
  END r0_rd_out[431]
  PIN r0_rd_out[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 435.825 767.060 435.895 767.200 ;
    END
  END r0_rd_out[432]
  PIN r0_rd_out[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 438.295 767.060 438.365 767.200 ;
    END
  END r0_rd_out[433]
  PIN r0_rd_out[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 440.765 767.060 440.835 767.200 ;
    END
  END r0_rd_out[434]
  PIN r0_rd_out[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 443.235 767.060 443.305 767.200 ;
    END
  END r0_rd_out[435]
  PIN r0_rd_out[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 445.705 767.060 445.775 767.200 ;
    END
  END r0_rd_out[436]
  PIN r0_rd_out[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 448.175 767.060 448.245 767.200 ;
    END
  END r0_rd_out[437]
  PIN r0_rd_out[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 450.645 767.060 450.715 767.200 ;
    END
  END r0_rd_out[438]
  PIN r0_rd_out[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 453.115 767.060 453.185 767.200 ;
    END
  END r0_rd_out[439]
  PIN r0_rd_out[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 455.585 767.060 455.655 767.200 ;
    END
  END r0_rd_out[440]
  PIN r0_rd_out[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 458.055 767.060 458.125 767.200 ;
    END
  END r0_rd_out[441]
  PIN r0_rd_out[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 460.525 767.060 460.595 767.200 ;
    END
  END r0_rd_out[442]
  PIN r0_rd_out[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 462.995 767.060 463.065 767.200 ;
    END
  END r0_rd_out[443]
  PIN r0_rd_out[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 465.465 767.060 465.535 767.200 ;
    END
  END r0_rd_out[444]
  PIN r0_rd_out[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 467.935 767.060 468.005 767.200 ;
    END
  END r0_rd_out[445]
  PIN r0_rd_out[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 470.405 767.060 470.475 767.200 ;
    END
  END r0_rd_out[446]
  PIN r0_rd_out[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 472.875 767.060 472.945 767.200 ;
    END
  END r0_rd_out[447]
  PIN r0_rd_out[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 475.345 767.060 475.415 767.200 ;
    END
  END r0_rd_out[448]
  PIN r0_rd_out[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 477.815 767.060 477.885 767.200 ;
    END
  END r0_rd_out[449]
  PIN r0_rd_out[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 480.285 767.060 480.355 767.200 ;
    END
  END r0_rd_out[450]
  PIN r0_rd_out[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 482.755 767.060 482.825 767.200 ;
    END
  END r0_rd_out[451]
  PIN r0_rd_out[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 485.225 767.060 485.295 767.200 ;
    END
  END r0_rd_out[452]
  PIN r0_rd_out[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 487.695 767.060 487.765 767.200 ;
    END
  END r0_rd_out[453]
  PIN r0_rd_out[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 490.165 767.060 490.235 767.200 ;
    END
  END r0_rd_out[454]
  PIN r0_rd_out[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 492.635 767.060 492.705 767.200 ;
    END
  END r0_rd_out[455]
  PIN r0_rd_out[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 495.105 767.060 495.175 767.200 ;
    END
  END r0_rd_out[456]
  PIN r0_rd_out[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 497.575 767.060 497.645 767.200 ;
    END
  END r0_rd_out[457]
  PIN r0_rd_out[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 500.045 767.060 500.115 767.200 ;
    END
  END r0_rd_out[458]
  PIN r0_rd_out[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 502.515 767.060 502.585 767.200 ;
    END
  END r0_rd_out[459]
  PIN r0_rd_out[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 504.985 767.060 505.055 767.200 ;
    END
  END r0_rd_out[460]
  PIN r0_rd_out[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 507.455 767.060 507.525 767.200 ;
    END
  END r0_rd_out[461]
  PIN r0_rd_out[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 509.925 767.060 509.995 767.200 ;
    END
  END r0_rd_out[462]
  PIN r0_rd_out[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 512.395 767.060 512.465 767.200 ;
    END
  END r0_rd_out[463]
  PIN r0_rd_out[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 514.865 767.060 514.935 767.200 ;
    END
  END r0_rd_out[464]
  PIN r0_rd_out[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 517.335 767.060 517.405 767.200 ;
    END
  END r0_rd_out[465]
  PIN r0_rd_out[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 519.805 767.060 519.875 767.200 ;
    END
  END r0_rd_out[466]
  PIN r0_rd_out[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 522.275 767.060 522.345 767.200 ;
    END
  END r0_rd_out[467]
  PIN r0_rd_out[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 524.745 767.060 524.815 767.200 ;
    END
  END r0_rd_out[468]
  PIN r0_rd_out[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 527.215 767.060 527.285 767.200 ;
    END
  END r0_rd_out[469]
  PIN r0_rd_out[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 529.685 767.060 529.755 767.200 ;
    END
  END r0_rd_out[470]
  PIN r0_rd_out[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 532.155 767.060 532.225 767.200 ;
    END
  END r0_rd_out[471]
  PIN r0_rd_out[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 534.625 767.060 534.695 767.200 ;
    END
  END r0_rd_out[472]
  PIN r0_rd_out[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 537.095 767.060 537.165 767.200 ;
    END
  END r0_rd_out[473]
  PIN r0_rd_out[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 539.565 767.060 539.635 767.200 ;
    END
  END r0_rd_out[474]
  PIN r0_rd_out[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 542.035 767.060 542.105 767.200 ;
    END
  END r0_rd_out[475]
  PIN r0_rd_out[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 544.505 767.060 544.575 767.200 ;
    END
  END r0_rd_out[476]
  PIN r0_rd_out[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 546.975 767.060 547.045 767.200 ;
    END
  END r0_rd_out[477]
  PIN r0_rd_out[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 549.445 767.060 549.515 767.200 ;
    END
  END r0_rd_out[478]
  PIN r0_rd_out[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 551.915 767.060 551.985 767.200 ;
    END
  END r0_rd_out[479]
  PIN r0_rd_out[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 554.385 767.060 554.455 767.200 ;
    END
  END r0_rd_out[480]
  PIN r0_rd_out[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 556.855 767.060 556.925 767.200 ;
    END
  END r0_rd_out[481]
  PIN r0_rd_out[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 559.325 767.060 559.395 767.200 ;
    END
  END r0_rd_out[482]
  PIN r0_rd_out[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 561.795 767.060 561.865 767.200 ;
    END
  END r0_rd_out[483]
  PIN r0_rd_out[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 564.265 767.060 564.335 767.200 ;
    END
  END r0_rd_out[484]
  PIN r0_rd_out[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 566.735 767.060 566.805 767.200 ;
    END
  END r0_rd_out[485]
  PIN r0_rd_out[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 569.205 767.060 569.275 767.200 ;
    END
  END r0_rd_out[486]
  PIN r0_rd_out[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 571.675 767.060 571.745 767.200 ;
    END
  END r0_rd_out[487]
  PIN r0_rd_out[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 574.145 767.060 574.215 767.200 ;
    END
  END r0_rd_out[488]
  PIN r0_rd_out[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 576.615 767.060 576.685 767.200 ;
    END
  END r0_rd_out[489]
  PIN r0_rd_out[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 579.085 767.060 579.155 767.200 ;
    END
  END r0_rd_out[490]
  PIN r0_rd_out[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 581.555 767.060 581.625 767.200 ;
    END
  END r0_rd_out[491]
  PIN r0_rd_out[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 584.025 767.060 584.095 767.200 ;
    END
  END r0_rd_out[492]
  PIN r0_rd_out[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 586.495 767.060 586.565 767.200 ;
    END
  END r0_rd_out[493]
  PIN r0_rd_out[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 588.965 767.060 589.035 767.200 ;
    END
  END r0_rd_out[494]
  PIN r0_rd_out[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 591.435 767.060 591.505 767.200 ;
    END
  END r0_rd_out[495]
  PIN r0_rd_out[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 593.905 767.060 593.975 767.200 ;
    END
  END r0_rd_out[496]
  PIN r0_rd_out[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 596.375 767.060 596.445 767.200 ;
    END
  END r0_rd_out[497]
  PIN r0_rd_out[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 598.845 767.060 598.915 767.200 ;
    END
  END r0_rd_out[498]
  PIN r0_rd_out[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 601.315 767.060 601.385 767.200 ;
    END
  END r0_rd_out[499]
  PIN r0_rd_out[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 603.785 767.060 603.855 767.200 ;
    END
  END r0_rd_out[500]
  PIN r0_rd_out[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 606.255 767.060 606.325 767.200 ;
    END
  END r0_rd_out[501]
  PIN r0_rd_out[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 608.725 767.060 608.795 767.200 ;
    END
  END r0_rd_out[502]
  PIN r0_rd_out[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 611.195 767.060 611.265 767.200 ;
    END
  END r0_rd_out[503]
  PIN r0_rd_out[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 613.665 767.060 613.735 767.200 ;
    END
  END r0_rd_out[504]
  PIN r0_rd_out[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 616.135 767.060 616.205 767.200 ;
    END
  END r0_rd_out[505]
  PIN r0_rd_out[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 618.605 767.060 618.675 767.200 ;
    END
  END r0_rd_out[506]
  PIN r0_rd_out[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 621.075 767.060 621.145 767.200 ;
    END
  END r0_rd_out[507]
  PIN r0_rd_out[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 623.545 767.060 623.615 767.200 ;
    END
  END r0_rd_out[508]
  PIN r0_rd_out[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 626.015 767.060 626.085 767.200 ;
    END
  END r0_rd_out[509]
  PIN r0_rd_out[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 628.485 767.060 628.555 767.200 ;
    END
  END r0_rd_out[510]
  PIN r0_rd_out[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 630.955 767.060 631.025 767.200 ;
    END
  END r0_rd_out[511]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.605 0.140 717.675 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.205 0.140 723.275 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 728.805 0.140 728.875 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 734.405 0.140 734.475 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 717.605 689.130 717.675 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 723.205 689.130 723.275 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 728.805 689.130 728.875 ;
    END
  END w0_addr_in[6]
  PIN w0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 734.405 689.130 734.475 ;
    END
  END w0_addr_in[7]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.005 0.140 740.075 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 745.605 0.140 745.675 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 751.205 0.140 751.275 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 756.805 0.140 756.875 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 740.005 689.130 740.075 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 745.605 689.130 745.675 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 751.205 689.130 751.275 ;
    END
  END r0_addr_in[6]
  PIN r0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 688.990 756.805 689.130 756.875 ;
    END
  END r0_addr_in[7]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 633.425 767.060 633.495 767.200 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 635.895 767.060 635.965 767.200 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 638.365 767.060 638.435 767.200 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 640.835 767.060 640.905 767.200 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 643.305 767.060 643.375 767.200 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 0.430 0.700 0.710 766.500 ;
      RECT 2.670 0.700 2.950 766.500 ;
      RECT 4.910 0.700 5.190 766.500 ;
      RECT 7.150 0.700 7.430 766.500 ;
      RECT 9.390 0.700 9.670 766.500 ;
      RECT 11.630 0.700 11.910 766.500 ;
      RECT 13.870 0.700 14.150 766.500 ;
      RECT 16.110 0.700 16.390 766.500 ;
      RECT 18.350 0.700 18.630 766.500 ;
      RECT 20.590 0.700 20.870 766.500 ;
      RECT 22.830 0.700 23.110 766.500 ;
      RECT 25.070 0.700 25.350 766.500 ;
      RECT 27.310 0.700 27.590 766.500 ;
      RECT 29.550 0.700 29.830 766.500 ;
      RECT 31.790 0.700 32.070 766.500 ;
      RECT 34.030 0.700 34.310 766.500 ;
      RECT 36.270 0.700 36.550 766.500 ;
      RECT 38.510 0.700 38.790 766.500 ;
      RECT 40.750 0.700 41.030 766.500 ;
      RECT 42.990 0.700 43.270 766.500 ;
      RECT 45.230 0.700 45.510 766.500 ;
      RECT 47.470 0.700 47.750 766.500 ;
      RECT 49.710 0.700 49.990 766.500 ;
      RECT 51.950 0.700 52.230 766.500 ;
      RECT 54.190 0.700 54.470 766.500 ;
      RECT 56.430 0.700 56.710 766.500 ;
      RECT 58.670 0.700 58.950 766.500 ;
      RECT 60.910 0.700 61.190 766.500 ;
      RECT 63.150 0.700 63.430 766.500 ;
      RECT 65.390 0.700 65.670 766.500 ;
      RECT 67.630 0.700 67.910 766.500 ;
      RECT 69.870 0.700 70.150 766.500 ;
      RECT 72.110 0.700 72.390 766.500 ;
      RECT 74.350 0.700 74.630 766.500 ;
      RECT 76.590 0.700 76.870 766.500 ;
      RECT 78.830 0.700 79.110 766.500 ;
      RECT 81.070 0.700 81.350 766.500 ;
      RECT 83.310 0.700 83.590 766.500 ;
      RECT 85.550 0.700 85.830 766.500 ;
      RECT 87.790 0.700 88.070 766.500 ;
      RECT 90.030 0.700 90.310 766.500 ;
      RECT 92.270 0.700 92.550 766.500 ;
      RECT 94.510 0.700 94.790 766.500 ;
      RECT 96.750 0.700 97.030 766.500 ;
      RECT 98.990 0.700 99.270 766.500 ;
      RECT 101.230 0.700 101.510 766.500 ;
      RECT 103.470 0.700 103.750 766.500 ;
      RECT 105.710 0.700 105.990 766.500 ;
      RECT 107.950 0.700 108.230 766.500 ;
      RECT 110.190 0.700 110.470 766.500 ;
      RECT 112.430 0.700 112.710 766.500 ;
      RECT 114.670 0.700 114.950 766.500 ;
      RECT 116.910 0.700 117.190 766.500 ;
      RECT 119.150 0.700 119.430 766.500 ;
      RECT 121.390 0.700 121.670 766.500 ;
      RECT 123.630 0.700 123.910 766.500 ;
      RECT 125.870 0.700 126.150 766.500 ;
      RECT 128.110 0.700 128.390 766.500 ;
      RECT 130.350 0.700 130.630 766.500 ;
      RECT 132.590 0.700 132.870 766.500 ;
      RECT 134.830 0.700 135.110 766.500 ;
      RECT 137.070 0.700 137.350 766.500 ;
      RECT 139.310 0.700 139.590 766.500 ;
      RECT 141.550 0.700 141.830 766.500 ;
      RECT 143.790 0.700 144.070 766.500 ;
      RECT 146.030 0.700 146.310 766.500 ;
      RECT 148.270 0.700 148.550 766.500 ;
      RECT 150.510 0.700 150.790 766.500 ;
      RECT 152.750 0.700 153.030 766.500 ;
      RECT 154.990 0.700 155.270 766.500 ;
      RECT 157.230 0.700 157.510 766.500 ;
      RECT 159.470 0.700 159.750 766.500 ;
      RECT 161.710 0.700 161.990 766.500 ;
      RECT 163.950 0.700 164.230 766.500 ;
      RECT 166.190 0.700 166.470 766.500 ;
      RECT 168.430 0.700 168.710 766.500 ;
      RECT 170.670 0.700 170.950 766.500 ;
      RECT 172.910 0.700 173.190 766.500 ;
      RECT 175.150 0.700 175.430 766.500 ;
      RECT 177.390 0.700 177.670 766.500 ;
      RECT 179.630 0.700 179.910 766.500 ;
      RECT 181.870 0.700 182.150 766.500 ;
      RECT 184.110 0.700 184.390 766.500 ;
      RECT 186.350 0.700 186.630 766.500 ;
      RECT 188.590 0.700 188.870 766.500 ;
      RECT 190.830 0.700 191.110 766.500 ;
      RECT 193.070 0.700 193.350 766.500 ;
      RECT 195.310 0.700 195.590 766.500 ;
      RECT 197.550 0.700 197.830 766.500 ;
      RECT 199.790 0.700 200.070 766.500 ;
      RECT 202.030 0.700 202.310 766.500 ;
      RECT 204.270 0.700 204.550 766.500 ;
      RECT 206.510 0.700 206.790 766.500 ;
      RECT 208.750 0.700 209.030 766.500 ;
      RECT 210.990 0.700 211.270 766.500 ;
      RECT 213.230 0.700 213.510 766.500 ;
      RECT 215.470 0.700 215.750 766.500 ;
      RECT 217.710 0.700 217.990 766.500 ;
      RECT 219.950 0.700 220.230 766.500 ;
      RECT 222.190 0.700 222.470 766.500 ;
      RECT 224.430 0.700 224.710 766.500 ;
      RECT 226.670 0.700 226.950 766.500 ;
      RECT 228.910 0.700 229.190 766.500 ;
      RECT 231.150 0.700 231.430 766.500 ;
      RECT 233.390 0.700 233.670 766.500 ;
      RECT 235.630 0.700 235.910 766.500 ;
      RECT 237.870 0.700 238.150 766.500 ;
      RECT 240.110 0.700 240.390 766.500 ;
      RECT 242.350 0.700 242.630 766.500 ;
      RECT 244.590 0.700 244.870 766.500 ;
      RECT 246.830 0.700 247.110 766.500 ;
      RECT 249.070 0.700 249.350 766.500 ;
      RECT 251.310 0.700 251.590 766.500 ;
      RECT 253.550 0.700 253.830 766.500 ;
      RECT 255.790 0.700 256.070 766.500 ;
      RECT 258.030 0.700 258.310 766.500 ;
      RECT 260.270 0.700 260.550 766.500 ;
      RECT 262.510 0.700 262.790 766.500 ;
      RECT 264.750 0.700 265.030 766.500 ;
      RECT 266.990 0.700 267.270 766.500 ;
      RECT 269.230 0.700 269.510 766.500 ;
      RECT 271.470 0.700 271.750 766.500 ;
      RECT 273.710 0.700 273.990 766.500 ;
      RECT 275.950 0.700 276.230 766.500 ;
      RECT 278.190 0.700 278.470 766.500 ;
      RECT 280.430 0.700 280.710 766.500 ;
      RECT 282.670 0.700 282.950 766.500 ;
      RECT 284.910 0.700 285.190 766.500 ;
      RECT 287.150 0.700 287.430 766.500 ;
      RECT 289.390 0.700 289.670 766.500 ;
      RECT 291.630 0.700 291.910 766.500 ;
      RECT 293.870 0.700 294.150 766.500 ;
      RECT 296.110 0.700 296.390 766.500 ;
      RECT 298.350 0.700 298.630 766.500 ;
      RECT 300.590 0.700 300.870 766.500 ;
      RECT 302.830 0.700 303.110 766.500 ;
      RECT 305.070 0.700 305.350 766.500 ;
      RECT 307.310 0.700 307.590 766.500 ;
      RECT 309.550 0.700 309.830 766.500 ;
      RECT 311.790 0.700 312.070 766.500 ;
      RECT 314.030 0.700 314.310 766.500 ;
      RECT 316.270 0.700 316.550 766.500 ;
      RECT 318.510 0.700 318.790 766.500 ;
      RECT 320.750 0.700 321.030 766.500 ;
      RECT 322.990 0.700 323.270 766.500 ;
      RECT 325.230 0.700 325.510 766.500 ;
      RECT 327.470 0.700 327.750 766.500 ;
      RECT 329.710 0.700 329.990 766.500 ;
      RECT 331.950 0.700 332.230 766.500 ;
      RECT 334.190 0.700 334.470 766.500 ;
      RECT 336.430 0.700 336.710 766.500 ;
      RECT 338.670 0.700 338.950 766.500 ;
      RECT 340.910 0.700 341.190 766.500 ;
      RECT 343.150 0.700 343.430 766.500 ;
      RECT 345.390 0.700 345.670 766.500 ;
      RECT 347.630 0.700 347.910 766.500 ;
      RECT 349.870 0.700 350.150 766.500 ;
      RECT 352.110 0.700 352.390 766.500 ;
      RECT 354.350 0.700 354.630 766.500 ;
      RECT 356.590 0.700 356.870 766.500 ;
      RECT 358.830 0.700 359.110 766.500 ;
      RECT 361.070 0.700 361.350 766.500 ;
      RECT 363.310 0.700 363.590 766.500 ;
      RECT 365.550 0.700 365.830 766.500 ;
      RECT 367.790 0.700 368.070 766.500 ;
      RECT 370.030 0.700 370.310 766.500 ;
      RECT 372.270 0.700 372.550 766.500 ;
      RECT 374.510 0.700 374.790 766.500 ;
      RECT 376.750 0.700 377.030 766.500 ;
      RECT 378.990 0.700 379.270 766.500 ;
      RECT 381.230 0.700 381.510 766.500 ;
      RECT 383.470 0.700 383.750 766.500 ;
      RECT 385.710 0.700 385.990 766.500 ;
      RECT 387.950 0.700 388.230 766.500 ;
      RECT 390.190 0.700 390.470 766.500 ;
      RECT 392.430 0.700 392.710 766.500 ;
      RECT 394.670 0.700 394.950 766.500 ;
      RECT 396.910 0.700 397.190 766.500 ;
      RECT 399.150 0.700 399.430 766.500 ;
      RECT 401.390 0.700 401.670 766.500 ;
      RECT 403.630 0.700 403.910 766.500 ;
      RECT 405.870 0.700 406.150 766.500 ;
      RECT 408.110 0.700 408.390 766.500 ;
      RECT 410.350 0.700 410.630 766.500 ;
      RECT 412.590 0.700 412.870 766.500 ;
      RECT 414.830 0.700 415.110 766.500 ;
      RECT 417.070 0.700 417.350 766.500 ;
      RECT 419.310 0.700 419.590 766.500 ;
      RECT 421.550 0.700 421.830 766.500 ;
      RECT 423.790 0.700 424.070 766.500 ;
      RECT 426.030 0.700 426.310 766.500 ;
      RECT 428.270 0.700 428.550 766.500 ;
      RECT 430.510 0.700 430.790 766.500 ;
      RECT 432.750 0.700 433.030 766.500 ;
      RECT 434.990 0.700 435.270 766.500 ;
      RECT 437.230 0.700 437.510 766.500 ;
      RECT 439.470 0.700 439.750 766.500 ;
      RECT 441.710 0.700 441.990 766.500 ;
      RECT 443.950 0.700 444.230 766.500 ;
      RECT 446.190 0.700 446.470 766.500 ;
      RECT 448.430 0.700 448.710 766.500 ;
      RECT 450.670 0.700 450.950 766.500 ;
      RECT 452.910 0.700 453.190 766.500 ;
      RECT 455.150 0.700 455.430 766.500 ;
      RECT 457.390 0.700 457.670 766.500 ;
      RECT 459.630 0.700 459.910 766.500 ;
      RECT 461.870 0.700 462.150 766.500 ;
      RECT 464.110 0.700 464.390 766.500 ;
      RECT 466.350 0.700 466.630 766.500 ;
      RECT 468.590 0.700 468.870 766.500 ;
      RECT 470.830 0.700 471.110 766.500 ;
      RECT 473.070 0.700 473.350 766.500 ;
      RECT 475.310 0.700 475.590 766.500 ;
      RECT 477.550 0.700 477.830 766.500 ;
      RECT 479.790 0.700 480.070 766.500 ;
      RECT 482.030 0.700 482.310 766.500 ;
      RECT 484.270 0.700 484.550 766.500 ;
      RECT 486.510 0.700 486.790 766.500 ;
      RECT 488.750 0.700 489.030 766.500 ;
      RECT 490.990 0.700 491.270 766.500 ;
      RECT 493.230 0.700 493.510 766.500 ;
      RECT 495.470 0.700 495.750 766.500 ;
      RECT 497.710 0.700 497.990 766.500 ;
      RECT 499.950 0.700 500.230 766.500 ;
      RECT 502.190 0.700 502.470 766.500 ;
      RECT 504.430 0.700 504.710 766.500 ;
      RECT 506.670 0.700 506.950 766.500 ;
      RECT 508.910 0.700 509.190 766.500 ;
      RECT 511.150 0.700 511.430 766.500 ;
      RECT 513.390 0.700 513.670 766.500 ;
      RECT 515.630 0.700 515.910 766.500 ;
      RECT 517.870 0.700 518.150 766.500 ;
      RECT 520.110 0.700 520.390 766.500 ;
      RECT 522.350 0.700 522.630 766.500 ;
      RECT 524.590 0.700 524.870 766.500 ;
      RECT 526.830 0.700 527.110 766.500 ;
      RECT 529.070 0.700 529.350 766.500 ;
      RECT 531.310 0.700 531.590 766.500 ;
      RECT 533.550 0.700 533.830 766.500 ;
      RECT 535.790 0.700 536.070 766.500 ;
      RECT 538.030 0.700 538.310 766.500 ;
      RECT 540.270 0.700 540.550 766.500 ;
      RECT 542.510 0.700 542.790 766.500 ;
      RECT 544.750 0.700 545.030 766.500 ;
      RECT 546.990 0.700 547.270 766.500 ;
      RECT 549.230 0.700 549.510 766.500 ;
      RECT 551.470 0.700 551.750 766.500 ;
      RECT 553.710 0.700 553.990 766.500 ;
      RECT 555.950 0.700 556.230 766.500 ;
      RECT 558.190 0.700 558.470 766.500 ;
      RECT 560.430 0.700 560.710 766.500 ;
      RECT 562.670 0.700 562.950 766.500 ;
      RECT 564.910 0.700 565.190 766.500 ;
      RECT 567.150 0.700 567.430 766.500 ;
      RECT 569.390 0.700 569.670 766.500 ;
      RECT 571.630 0.700 571.910 766.500 ;
      RECT 573.870 0.700 574.150 766.500 ;
      RECT 576.110 0.700 576.390 766.500 ;
      RECT 578.350 0.700 578.630 766.500 ;
      RECT 580.590 0.700 580.870 766.500 ;
      RECT 582.830 0.700 583.110 766.500 ;
      RECT 585.070 0.700 585.350 766.500 ;
      RECT 587.310 0.700 587.590 766.500 ;
      RECT 589.550 0.700 589.830 766.500 ;
      RECT 591.790 0.700 592.070 766.500 ;
      RECT 594.030 0.700 594.310 766.500 ;
      RECT 596.270 0.700 596.550 766.500 ;
      RECT 598.510 0.700 598.790 766.500 ;
      RECT 600.750 0.700 601.030 766.500 ;
      RECT 602.990 0.700 603.270 766.500 ;
      RECT 605.230 0.700 605.510 766.500 ;
      RECT 607.470 0.700 607.750 766.500 ;
      RECT 609.710 0.700 609.990 766.500 ;
      RECT 611.950 0.700 612.230 766.500 ;
      RECT 614.190 0.700 614.470 766.500 ;
      RECT 616.430 0.700 616.710 766.500 ;
      RECT 618.670 0.700 618.950 766.500 ;
      RECT 620.910 0.700 621.190 766.500 ;
      RECT 623.150 0.700 623.430 766.500 ;
      RECT 625.390 0.700 625.670 766.500 ;
      RECT 627.630 0.700 627.910 766.500 ;
      RECT 629.870 0.700 630.150 766.500 ;
      RECT 632.110 0.700 632.390 766.500 ;
      RECT 634.350 0.700 634.630 766.500 ;
      RECT 636.590 0.700 636.870 766.500 ;
      RECT 638.830 0.700 639.110 766.500 ;
      RECT 641.070 0.700 641.350 766.500 ;
      RECT 643.310 0.700 643.590 766.500 ;
      RECT 645.550 0.700 645.830 766.500 ;
      RECT 647.790 0.700 648.070 766.500 ;
      RECT 650.030 0.700 650.310 766.500 ;
      RECT 652.270 0.700 652.550 766.500 ;
      RECT 654.510 0.700 654.790 766.500 ;
      RECT 656.750 0.700 657.030 766.500 ;
      RECT 658.990 0.700 659.270 766.500 ;
      RECT 661.230 0.700 661.510 766.500 ;
      RECT 663.470 0.700 663.750 766.500 ;
      RECT 665.710 0.700 665.990 766.500 ;
      RECT 667.950 0.700 668.230 766.500 ;
      RECT 670.190 0.700 670.470 766.500 ;
      RECT 672.430 0.700 672.710 766.500 ;
      RECT 674.670 0.700 674.950 766.500 ;
      RECT 676.910 0.700 677.190 766.500 ;
      RECT 679.150 0.700 679.430 766.500 ;
      RECT 681.390 0.700 681.670 766.500 ;
      RECT 683.630 0.700 683.910 766.500 ;
      RECT 685.870 0.700 686.150 766.500 ;
      RECT 688.110 0.700 688.390 766.500 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 0.430 0.700 0.710 766.500 ;
      RECT 2.670 0.700 2.950 766.500 ;
      RECT 4.910 0.700 5.190 766.500 ;
      RECT 7.150 0.700 7.430 766.500 ;
      RECT 9.390 0.700 9.670 766.500 ;
      RECT 11.630 0.700 11.910 766.500 ;
      RECT 13.870 0.700 14.150 766.500 ;
      RECT 16.110 0.700 16.390 766.500 ;
      RECT 18.350 0.700 18.630 766.500 ;
      RECT 20.590 0.700 20.870 766.500 ;
      RECT 22.830 0.700 23.110 766.500 ;
      RECT 25.070 0.700 25.350 766.500 ;
      RECT 27.310 0.700 27.590 766.500 ;
      RECT 29.550 0.700 29.830 766.500 ;
      RECT 31.790 0.700 32.070 766.500 ;
      RECT 34.030 0.700 34.310 766.500 ;
      RECT 36.270 0.700 36.550 766.500 ;
      RECT 38.510 0.700 38.790 766.500 ;
      RECT 40.750 0.700 41.030 766.500 ;
      RECT 42.990 0.700 43.270 766.500 ;
      RECT 45.230 0.700 45.510 766.500 ;
      RECT 47.470 0.700 47.750 766.500 ;
      RECT 49.710 0.700 49.990 766.500 ;
      RECT 51.950 0.700 52.230 766.500 ;
      RECT 54.190 0.700 54.470 766.500 ;
      RECT 56.430 0.700 56.710 766.500 ;
      RECT 58.670 0.700 58.950 766.500 ;
      RECT 60.910 0.700 61.190 766.500 ;
      RECT 63.150 0.700 63.430 766.500 ;
      RECT 65.390 0.700 65.670 766.500 ;
      RECT 67.630 0.700 67.910 766.500 ;
      RECT 69.870 0.700 70.150 766.500 ;
      RECT 72.110 0.700 72.390 766.500 ;
      RECT 74.350 0.700 74.630 766.500 ;
      RECT 76.590 0.700 76.870 766.500 ;
      RECT 78.830 0.700 79.110 766.500 ;
      RECT 81.070 0.700 81.350 766.500 ;
      RECT 83.310 0.700 83.590 766.500 ;
      RECT 85.550 0.700 85.830 766.500 ;
      RECT 87.790 0.700 88.070 766.500 ;
      RECT 90.030 0.700 90.310 766.500 ;
      RECT 92.270 0.700 92.550 766.500 ;
      RECT 94.510 0.700 94.790 766.500 ;
      RECT 96.750 0.700 97.030 766.500 ;
      RECT 98.990 0.700 99.270 766.500 ;
      RECT 101.230 0.700 101.510 766.500 ;
      RECT 103.470 0.700 103.750 766.500 ;
      RECT 105.710 0.700 105.990 766.500 ;
      RECT 107.950 0.700 108.230 766.500 ;
      RECT 110.190 0.700 110.470 766.500 ;
      RECT 112.430 0.700 112.710 766.500 ;
      RECT 114.670 0.700 114.950 766.500 ;
      RECT 116.910 0.700 117.190 766.500 ;
      RECT 119.150 0.700 119.430 766.500 ;
      RECT 121.390 0.700 121.670 766.500 ;
      RECT 123.630 0.700 123.910 766.500 ;
      RECT 125.870 0.700 126.150 766.500 ;
      RECT 128.110 0.700 128.390 766.500 ;
      RECT 130.350 0.700 130.630 766.500 ;
      RECT 132.590 0.700 132.870 766.500 ;
      RECT 134.830 0.700 135.110 766.500 ;
      RECT 137.070 0.700 137.350 766.500 ;
      RECT 139.310 0.700 139.590 766.500 ;
      RECT 141.550 0.700 141.830 766.500 ;
      RECT 143.790 0.700 144.070 766.500 ;
      RECT 146.030 0.700 146.310 766.500 ;
      RECT 148.270 0.700 148.550 766.500 ;
      RECT 150.510 0.700 150.790 766.500 ;
      RECT 152.750 0.700 153.030 766.500 ;
      RECT 154.990 0.700 155.270 766.500 ;
      RECT 157.230 0.700 157.510 766.500 ;
      RECT 159.470 0.700 159.750 766.500 ;
      RECT 161.710 0.700 161.990 766.500 ;
      RECT 163.950 0.700 164.230 766.500 ;
      RECT 166.190 0.700 166.470 766.500 ;
      RECT 168.430 0.700 168.710 766.500 ;
      RECT 170.670 0.700 170.950 766.500 ;
      RECT 172.910 0.700 173.190 766.500 ;
      RECT 175.150 0.700 175.430 766.500 ;
      RECT 177.390 0.700 177.670 766.500 ;
      RECT 179.630 0.700 179.910 766.500 ;
      RECT 181.870 0.700 182.150 766.500 ;
      RECT 184.110 0.700 184.390 766.500 ;
      RECT 186.350 0.700 186.630 766.500 ;
      RECT 188.590 0.700 188.870 766.500 ;
      RECT 190.830 0.700 191.110 766.500 ;
      RECT 193.070 0.700 193.350 766.500 ;
      RECT 195.310 0.700 195.590 766.500 ;
      RECT 197.550 0.700 197.830 766.500 ;
      RECT 199.790 0.700 200.070 766.500 ;
      RECT 202.030 0.700 202.310 766.500 ;
      RECT 204.270 0.700 204.550 766.500 ;
      RECT 206.510 0.700 206.790 766.500 ;
      RECT 208.750 0.700 209.030 766.500 ;
      RECT 210.990 0.700 211.270 766.500 ;
      RECT 213.230 0.700 213.510 766.500 ;
      RECT 215.470 0.700 215.750 766.500 ;
      RECT 217.710 0.700 217.990 766.500 ;
      RECT 219.950 0.700 220.230 766.500 ;
      RECT 222.190 0.700 222.470 766.500 ;
      RECT 224.430 0.700 224.710 766.500 ;
      RECT 226.670 0.700 226.950 766.500 ;
      RECT 228.910 0.700 229.190 766.500 ;
      RECT 231.150 0.700 231.430 766.500 ;
      RECT 233.390 0.700 233.670 766.500 ;
      RECT 235.630 0.700 235.910 766.500 ;
      RECT 237.870 0.700 238.150 766.500 ;
      RECT 240.110 0.700 240.390 766.500 ;
      RECT 242.350 0.700 242.630 766.500 ;
      RECT 244.590 0.700 244.870 766.500 ;
      RECT 246.830 0.700 247.110 766.500 ;
      RECT 249.070 0.700 249.350 766.500 ;
      RECT 251.310 0.700 251.590 766.500 ;
      RECT 253.550 0.700 253.830 766.500 ;
      RECT 255.790 0.700 256.070 766.500 ;
      RECT 258.030 0.700 258.310 766.500 ;
      RECT 260.270 0.700 260.550 766.500 ;
      RECT 262.510 0.700 262.790 766.500 ;
      RECT 264.750 0.700 265.030 766.500 ;
      RECT 266.990 0.700 267.270 766.500 ;
      RECT 269.230 0.700 269.510 766.500 ;
      RECT 271.470 0.700 271.750 766.500 ;
      RECT 273.710 0.700 273.990 766.500 ;
      RECT 275.950 0.700 276.230 766.500 ;
      RECT 278.190 0.700 278.470 766.500 ;
      RECT 280.430 0.700 280.710 766.500 ;
      RECT 282.670 0.700 282.950 766.500 ;
      RECT 284.910 0.700 285.190 766.500 ;
      RECT 287.150 0.700 287.430 766.500 ;
      RECT 289.390 0.700 289.670 766.500 ;
      RECT 291.630 0.700 291.910 766.500 ;
      RECT 293.870 0.700 294.150 766.500 ;
      RECT 296.110 0.700 296.390 766.500 ;
      RECT 298.350 0.700 298.630 766.500 ;
      RECT 300.590 0.700 300.870 766.500 ;
      RECT 302.830 0.700 303.110 766.500 ;
      RECT 305.070 0.700 305.350 766.500 ;
      RECT 307.310 0.700 307.590 766.500 ;
      RECT 309.550 0.700 309.830 766.500 ;
      RECT 311.790 0.700 312.070 766.500 ;
      RECT 314.030 0.700 314.310 766.500 ;
      RECT 316.270 0.700 316.550 766.500 ;
      RECT 318.510 0.700 318.790 766.500 ;
      RECT 320.750 0.700 321.030 766.500 ;
      RECT 322.990 0.700 323.270 766.500 ;
      RECT 325.230 0.700 325.510 766.500 ;
      RECT 327.470 0.700 327.750 766.500 ;
      RECT 329.710 0.700 329.990 766.500 ;
      RECT 331.950 0.700 332.230 766.500 ;
      RECT 334.190 0.700 334.470 766.500 ;
      RECT 336.430 0.700 336.710 766.500 ;
      RECT 338.670 0.700 338.950 766.500 ;
      RECT 340.910 0.700 341.190 766.500 ;
      RECT 343.150 0.700 343.430 766.500 ;
      RECT 345.390 0.700 345.670 766.500 ;
      RECT 347.630 0.700 347.910 766.500 ;
      RECT 349.870 0.700 350.150 766.500 ;
      RECT 352.110 0.700 352.390 766.500 ;
      RECT 354.350 0.700 354.630 766.500 ;
      RECT 356.590 0.700 356.870 766.500 ;
      RECT 358.830 0.700 359.110 766.500 ;
      RECT 361.070 0.700 361.350 766.500 ;
      RECT 363.310 0.700 363.590 766.500 ;
      RECT 365.550 0.700 365.830 766.500 ;
      RECT 367.790 0.700 368.070 766.500 ;
      RECT 370.030 0.700 370.310 766.500 ;
      RECT 372.270 0.700 372.550 766.500 ;
      RECT 374.510 0.700 374.790 766.500 ;
      RECT 376.750 0.700 377.030 766.500 ;
      RECT 378.990 0.700 379.270 766.500 ;
      RECT 381.230 0.700 381.510 766.500 ;
      RECT 383.470 0.700 383.750 766.500 ;
      RECT 385.710 0.700 385.990 766.500 ;
      RECT 387.950 0.700 388.230 766.500 ;
      RECT 390.190 0.700 390.470 766.500 ;
      RECT 392.430 0.700 392.710 766.500 ;
      RECT 394.670 0.700 394.950 766.500 ;
      RECT 396.910 0.700 397.190 766.500 ;
      RECT 399.150 0.700 399.430 766.500 ;
      RECT 401.390 0.700 401.670 766.500 ;
      RECT 403.630 0.700 403.910 766.500 ;
      RECT 405.870 0.700 406.150 766.500 ;
      RECT 408.110 0.700 408.390 766.500 ;
      RECT 410.350 0.700 410.630 766.500 ;
      RECT 412.590 0.700 412.870 766.500 ;
      RECT 414.830 0.700 415.110 766.500 ;
      RECT 417.070 0.700 417.350 766.500 ;
      RECT 419.310 0.700 419.590 766.500 ;
      RECT 421.550 0.700 421.830 766.500 ;
      RECT 423.790 0.700 424.070 766.500 ;
      RECT 426.030 0.700 426.310 766.500 ;
      RECT 428.270 0.700 428.550 766.500 ;
      RECT 430.510 0.700 430.790 766.500 ;
      RECT 432.750 0.700 433.030 766.500 ;
      RECT 434.990 0.700 435.270 766.500 ;
      RECT 437.230 0.700 437.510 766.500 ;
      RECT 439.470 0.700 439.750 766.500 ;
      RECT 441.710 0.700 441.990 766.500 ;
      RECT 443.950 0.700 444.230 766.500 ;
      RECT 446.190 0.700 446.470 766.500 ;
      RECT 448.430 0.700 448.710 766.500 ;
      RECT 450.670 0.700 450.950 766.500 ;
      RECT 452.910 0.700 453.190 766.500 ;
      RECT 455.150 0.700 455.430 766.500 ;
      RECT 457.390 0.700 457.670 766.500 ;
      RECT 459.630 0.700 459.910 766.500 ;
      RECT 461.870 0.700 462.150 766.500 ;
      RECT 464.110 0.700 464.390 766.500 ;
      RECT 466.350 0.700 466.630 766.500 ;
      RECT 468.590 0.700 468.870 766.500 ;
      RECT 470.830 0.700 471.110 766.500 ;
      RECT 473.070 0.700 473.350 766.500 ;
      RECT 475.310 0.700 475.590 766.500 ;
      RECT 477.550 0.700 477.830 766.500 ;
      RECT 479.790 0.700 480.070 766.500 ;
      RECT 482.030 0.700 482.310 766.500 ;
      RECT 484.270 0.700 484.550 766.500 ;
      RECT 486.510 0.700 486.790 766.500 ;
      RECT 488.750 0.700 489.030 766.500 ;
      RECT 490.990 0.700 491.270 766.500 ;
      RECT 493.230 0.700 493.510 766.500 ;
      RECT 495.470 0.700 495.750 766.500 ;
      RECT 497.710 0.700 497.990 766.500 ;
      RECT 499.950 0.700 500.230 766.500 ;
      RECT 502.190 0.700 502.470 766.500 ;
      RECT 504.430 0.700 504.710 766.500 ;
      RECT 506.670 0.700 506.950 766.500 ;
      RECT 508.910 0.700 509.190 766.500 ;
      RECT 511.150 0.700 511.430 766.500 ;
      RECT 513.390 0.700 513.670 766.500 ;
      RECT 515.630 0.700 515.910 766.500 ;
      RECT 517.870 0.700 518.150 766.500 ;
      RECT 520.110 0.700 520.390 766.500 ;
      RECT 522.350 0.700 522.630 766.500 ;
      RECT 524.590 0.700 524.870 766.500 ;
      RECT 526.830 0.700 527.110 766.500 ;
      RECT 529.070 0.700 529.350 766.500 ;
      RECT 531.310 0.700 531.590 766.500 ;
      RECT 533.550 0.700 533.830 766.500 ;
      RECT 535.790 0.700 536.070 766.500 ;
      RECT 538.030 0.700 538.310 766.500 ;
      RECT 540.270 0.700 540.550 766.500 ;
      RECT 542.510 0.700 542.790 766.500 ;
      RECT 544.750 0.700 545.030 766.500 ;
      RECT 546.990 0.700 547.270 766.500 ;
      RECT 549.230 0.700 549.510 766.500 ;
      RECT 551.470 0.700 551.750 766.500 ;
      RECT 553.710 0.700 553.990 766.500 ;
      RECT 555.950 0.700 556.230 766.500 ;
      RECT 558.190 0.700 558.470 766.500 ;
      RECT 560.430 0.700 560.710 766.500 ;
      RECT 562.670 0.700 562.950 766.500 ;
      RECT 564.910 0.700 565.190 766.500 ;
      RECT 567.150 0.700 567.430 766.500 ;
      RECT 569.390 0.700 569.670 766.500 ;
      RECT 571.630 0.700 571.910 766.500 ;
      RECT 573.870 0.700 574.150 766.500 ;
      RECT 576.110 0.700 576.390 766.500 ;
      RECT 578.350 0.700 578.630 766.500 ;
      RECT 580.590 0.700 580.870 766.500 ;
      RECT 582.830 0.700 583.110 766.500 ;
      RECT 585.070 0.700 585.350 766.500 ;
      RECT 587.310 0.700 587.590 766.500 ;
      RECT 589.550 0.700 589.830 766.500 ;
      RECT 591.790 0.700 592.070 766.500 ;
      RECT 594.030 0.700 594.310 766.500 ;
      RECT 596.270 0.700 596.550 766.500 ;
      RECT 598.510 0.700 598.790 766.500 ;
      RECT 600.750 0.700 601.030 766.500 ;
      RECT 602.990 0.700 603.270 766.500 ;
      RECT 605.230 0.700 605.510 766.500 ;
      RECT 607.470 0.700 607.750 766.500 ;
      RECT 609.710 0.700 609.990 766.500 ;
      RECT 611.950 0.700 612.230 766.500 ;
      RECT 614.190 0.700 614.470 766.500 ;
      RECT 616.430 0.700 616.710 766.500 ;
      RECT 618.670 0.700 618.950 766.500 ;
      RECT 620.910 0.700 621.190 766.500 ;
      RECT 623.150 0.700 623.430 766.500 ;
      RECT 625.390 0.700 625.670 766.500 ;
      RECT 627.630 0.700 627.910 766.500 ;
      RECT 629.870 0.700 630.150 766.500 ;
      RECT 632.110 0.700 632.390 766.500 ;
      RECT 634.350 0.700 634.630 766.500 ;
      RECT 636.590 0.700 636.870 766.500 ;
      RECT 638.830 0.700 639.110 766.500 ;
      RECT 641.070 0.700 641.350 766.500 ;
      RECT 643.310 0.700 643.590 766.500 ;
      RECT 645.550 0.700 645.830 766.500 ;
      RECT 647.790 0.700 648.070 766.500 ;
      RECT 650.030 0.700 650.310 766.500 ;
      RECT 652.270 0.700 652.550 766.500 ;
      RECT 654.510 0.700 654.790 766.500 ;
      RECT 656.750 0.700 657.030 766.500 ;
      RECT 658.990 0.700 659.270 766.500 ;
      RECT 661.230 0.700 661.510 766.500 ;
      RECT 663.470 0.700 663.750 766.500 ;
      RECT 665.710 0.700 665.990 766.500 ;
      RECT 667.950 0.700 668.230 766.500 ;
      RECT 670.190 0.700 670.470 766.500 ;
      RECT 672.430 0.700 672.710 766.500 ;
      RECT 674.670 0.700 674.950 766.500 ;
      RECT 676.910 0.700 677.190 766.500 ;
      RECT 679.150 0.700 679.430 766.500 ;
      RECT 681.390 0.700 681.670 766.500 ;
      RECT 683.630 0.700 683.910 766.500 ;
      RECT 685.870 0.700 686.150 766.500 ;
      RECT 688.110 0.700 688.390 766.500 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 689.130 767.200 ;
    LAYER metal2 ;
    RECT 0 0 689.130 767.200 ;
    LAYER metal3 ;
    RECT 0 0 689.130 767.200 ;
    LAYER metal4 ;
    RECT 0 0 689.130 767.200 ;
    LAYER OVERLAP ;
    RECT 0 0 689.130 767.200 ;
  END
END fakeram_512x256_1r1w

END LIBRARY
