VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_20x64_1r1w
  FOREIGN fakeram_20x64_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 76.950 BY 63.000 ;
  CLASS BLOCK ;
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 0.805 0.140 0.875 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.140 6.335 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.140 11.795 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.140 17.255 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.140 22.715 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 76.810 0.805 76.950 0.875 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 76.810 6.265 76.950 6.335 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 76.810 11.725 76.950 11.795 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 76.810 17.185 76.950 17.255 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 76.810 22.645 76.950 22.715 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1.105 0.000 1.175 0.140 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 4.715 0.000 4.785 0.140 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 8.325 0.000 8.395 0.140 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 11.935 0.000 12.005 0.140 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 15.545 0.000 15.615 0.140 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 19.155 0.000 19.225 0.140 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 22.765 0.000 22.835 0.140 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 26.375 0.000 26.445 0.140 ;
    END
  END w0_wd_in[17]
  PIN w0_wd_in[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 29.985 0.000 30.055 0.140 ;
    END
  END w0_wd_in[18]
  PIN w0_wd_in[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 33.595 0.000 33.665 0.140 ;
    END
  END w0_wd_in[19]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 37.205 0.000 37.275 0.140 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 40.815 0.000 40.885 0.140 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 44.425 0.000 44.495 0.140 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 48.035 0.000 48.105 0.140 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 51.645 0.000 51.715 0.140 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 55.255 0.000 55.325 0.140 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 58.865 0.000 58.935 0.140 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 62.475 0.000 62.545 0.140 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 66.085 0.000 66.155 0.140 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 69.695 0.000 69.765 0.140 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1.105 62.860 1.175 63.000 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 6.045 62.860 6.115 63.000 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 10.985 62.860 11.055 63.000 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 15.925 62.860 15.995 63.000 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 20.865 62.860 20.935 63.000 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 25.805 62.860 25.875 63.000 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 30.745 62.860 30.815 63.000 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 35.685 62.860 35.755 63.000 ;
    END
  END r0_rd_out[17]
  PIN r0_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 40.625 62.860 40.695 63.000 ;
    END
  END r0_rd_out[18]
  PIN r0_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 45.565 62.860 45.635 63.000 ;
    END
  END r0_rd_out[19]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.105 0.140 28.175 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.140 33.635 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.140 39.095 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 76.810 28.105 76.950 28.175 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 76.810 33.565 76.950 33.635 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 76.810 39.025 76.950 39.095 ;
    END
  END w0_addr_in[5]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.140 44.555 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.140 50.015 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.140 55.475 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 76.810 44.485 76.950 44.555 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 76.810 49.945 76.950 50.015 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 76.810 55.405 76.950 55.475 ;
    END
  END r0_addr_in[5]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 50.505 62.860 50.575 63.000 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 55.445 62.860 55.515 63.000 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 60.385 62.860 60.455 63.000 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 65.325 62.860 65.395 63.000 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 70.265 62.860 70.335 63.000 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 0.430 0.700 0.710 62.300 ;
      RECT 2.670 0.700 2.950 62.300 ;
      RECT 4.910 0.700 5.190 62.300 ;
      RECT 7.150 0.700 7.430 62.300 ;
      RECT 9.390 0.700 9.670 62.300 ;
      RECT 11.630 0.700 11.910 62.300 ;
      RECT 13.870 0.700 14.150 62.300 ;
      RECT 16.110 0.700 16.390 62.300 ;
      RECT 18.350 0.700 18.630 62.300 ;
      RECT 20.590 0.700 20.870 62.300 ;
      RECT 22.830 0.700 23.110 62.300 ;
      RECT 25.070 0.700 25.350 62.300 ;
      RECT 27.310 0.700 27.590 62.300 ;
      RECT 29.550 0.700 29.830 62.300 ;
      RECT 31.790 0.700 32.070 62.300 ;
      RECT 34.030 0.700 34.310 62.300 ;
      RECT 36.270 0.700 36.550 62.300 ;
      RECT 38.510 0.700 38.790 62.300 ;
      RECT 40.750 0.700 41.030 62.300 ;
      RECT 42.990 0.700 43.270 62.300 ;
      RECT 45.230 0.700 45.510 62.300 ;
      RECT 47.470 0.700 47.750 62.300 ;
      RECT 49.710 0.700 49.990 62.300 ;
      RECT 51.950 0.700 52.230 62.300 ;
      RECT 54.190 0.700 54.470 62.300 ;
      RECT 56.430 0.700 56.710 62.300 ;
      RECT 58.670 0.700 58.950 62.300 ;
      RECT 60.910 0.700 61.190 62.300 ;
      RECT 63.150 0.700 63.430 62.300 ;
      RECT 65.390 0.700 65.670 62.300 ;
      RECT 67.630 0.700 67.910 62.300 ;
      RECT 69.870 0.700 70.150 62.300 ;
      RECT 72.110 0.700 72.390 62.300 ;
      RECT 74.350 0.700 74.630 62.300 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 0.430 0.700 0.710 62.300 ;
      RECT 2.670 0.700 2.950 62.300 ;
      RECT 4.910 0.700 5.190 62.300 ;
      RECT 7.150 0.700 7.430 62.300 ;
      RECT 9.390 0.700 9.670 62.300 ;
      RECT 11.630 0.700 11.910 62.300 ;
      RECT 13.870 0.700 14.150 62.300 ;
      RECT 16.110 0.700 16.390 62.300 ;
      RECT 18.350 0.700 18.630 62.300 ;
      RECT 20.590 0.700 20.870 62.300 ;
      RECT 22.830 0.700 23.110 62.300 ;
      RECT 25.070 0.700 25.350 62.300 ;
      RECT 27.310 0.700 27.590 62.300 ;
      RECT 29.550 0.700 29.830 62.300 ;
      RECT 31.790 0.700 32.070 62.300 ;
      RECT 34.030 0.700 34.310 62.300 ;
      RECT 36.270 0.700 36.550 62.300 ;
      RECT 38.510 0.700 38.790 62.300 ;
      RECT 40.750 0.700 41.030 62.300 ;
      RECT 42.990 0.700 43.270 62.300 ;
      RECT 45.230 0.700 45.510 62.300 ;
      RECT 47.470 0.700 47.750 62.300 ;
      RECT 49.710 0.700 49.990 62.300 ;
      RECT 51.950 0.700 52.230 62.300 ;
      RECT 54.190 0.700 54.470 62.300 ;
      RECT 56.430 0.700 56.710 62.300 ;
      RECT 58.670 0.700 58.950 62.300 ;
      RECT 60.910 0.700 61.190 62.300 ;
      RECT 63.150 0.700 63.430 62.300 ;
      RECT 65.390 0.700 65.670 62.300 ;
      RECT 67.630 0.700 67.910 62.300 ;
      RECT 69.870 0.700 70.150 62.300 ;
      RECT 72.110 0.700 72.390 62.300 ;
      RECT 74.350 0.700 74.630 62.300 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 76.950 63.000 ;
    LAYER metal2 ;
    RECT 0 0 76.950 63.000 ;
    LAYER metal3 ;
    RECT 0 0 76.950 63.000 ;
    LAYER metal4 ;
    RECT 0 0 76.950 63.000 ;
    LAYER OVERLAP ;
    RECT 0 0 76.950 63.000 ;
  END
END fakeram_20x64_1r1w

END LIBRARY
