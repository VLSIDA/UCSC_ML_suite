VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_20x64_2r1w
  FOREIGN fakeram_20x64_2r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 477.940 BY 190.400 ;
  CLASS BLOCK ;
  PIN w0_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 6.650 0.800 6.950 ;
    END
  END w0_mask_in[0]
  PIN w0_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 10.730 0.800 11.030 ;
    END
  END w0_mask_in[1]
  PIN w0_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.810 0.800 15.110 ;
    END
  END w0_mask_in[2]
  PIN w0_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 18.890 0.800 19.190 ;
    END
  END w0_mask_in[3]
  PIN w0_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.970 0.800 23.270 ;
    END
  END w0_mask_in[4]
  PIN w0_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 27.050 0.800 27.350 ;
    END
  END w0_mask_in[5]
  PIN w0_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.130 0.800 31.430 ;
    END
  END w0_mask_in[6]
  PIN w0_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 35.210 0.800 35.510 ;
    END
  END w0_mask_in[7]
  PIN w0_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.290 0.800 39.590 ;
    END
  END w0_mask_in[8]
  PIN w0_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 43.370 0.800 43.670 ;
    END
  END w0_mask_in[9]
  PIN w0_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 47.450 0.800 47.750 ;
    END
  END w0_mask_in[10]
  PIN w0_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 51.530 0.800 51.830 ;
    END
  END w0_mask_in[11]
  PIN w0_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.610 0.800 55.910 ;
    END
  END w0_mask_in[12]
  PIN w0_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 59.690 0.800 59.990 ;
    END
  END w0_mask_in[13]
  PIN w0_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 63.770 0.800 64.070 ;
    END
  END w0_mask_in[14]
  PIN w0_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.850 0.800 68.150 ;
    END
  END w0_mask_in[15]
  PIN w0_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.930 0.800 72.230 ;
    END
  END w0_mask_in[16]
  PIN w0_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.010 0.800 76.310 ;
    END
  END w0_mask_in[17]
  PIN w0_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 80.090 0.800 80.390 ;
    END
  END w0_mask_in[18]
  PIN w0_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 84.170 0.800 84.470 ;
    END
  END w0_mask_in[19]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 90.970 0.800 91.270 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 95.050 0.800 95.350 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 99.130 0.800 99.430 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 103.210 0.800 103.510 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 107.290 0.800 107.590 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 111.370 0.800 111.670 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 115.450 0.800 115.750 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 119.530 0.800 119.830 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 123.610 0.800 123.910 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 127.690 0.800 127.990 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 131.770 0.800 132.070 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 135.850 0.800 136.150 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.930 0.800 140.230 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 144.010 0.800 144.310 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 148.090 0.800 148.390 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 152.170 0.800 152.470 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 156.250 0.800 156.550 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 160.330 0.800 160.630 ;
    END
  END w0_wd_in[17]
  PIN w0_wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 164.410 0.800 164.710 ;
    END
  END w0_wd_in[18]
  PIN w0_wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 168.490 0.800 168.790 ;
    END
  END w0_wd_in[19]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 0.000 4.670 0.350 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 16.030 0.000 16.170 0.350 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 27.530 0.000 27.670 0.350 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 39.030 0.000 39.170 0.350 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 50.530 0.000 50.670 0.350 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 62.030 0.000 62.170 0.350 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 73.530 0.000 73.670 0.350 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 85.030 0.000 85.170 0.350 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 96.530 0.000 96.670 0.350 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 108.030 0.000 108.170 0.350 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 119.530 0.000 119.670 0.350 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 131.030 0.000 131.170 0.350 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 142.530 0.000 142.670 0.350 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 154.030 0.000 154.170 0.350 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 165.530 0.000 165.670 0.350 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 177.030 0.000 177.170 0.350 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 188.530 0.000 188.670 0.350 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 200.030 0.000 200.170 0.350 ;
    END
  END r0_rd_out[17]
  PIN r0_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 211.530 0.000 211.670 0.350 ;
    END
  END r0_rd_out[18]
  PIN r0_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 223.030 0.000 223.170 0.350 ;
    END
  END r0_rd_out[19]
  PIN r1_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 227.170 0.000 227.310 0.350 ;
    END
  END r1_rd_out[0]
  PIN r1_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 238.670 0.000 238.810 0.350 ;
    END
  END r1_rd_out[1]
  PIN r1_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 250.170 0.000 250.310 0.350 ;
    END
  END r1_rd_out[2]
  PIN r1_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 261.670 0.000 261.810 0.350 ;
    END
  END r1_rd_out[3]
  PIN r1_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 273.170 0.000 273.310 0.350 ;
    END
  END r1_rd_out[4]
  PIN r1_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 284.670 0.000 284.810 0.350 ;
    END
  END r1_rd_out[5]
  PIN r1_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 296.170 0.000 296.310 0.350 ;
    END
  END r1_rd_out[6]
  PIN r1_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 307.670 0.000 307.810 0.350 ;
    END
  END r1_rd_out[7]
  PIN r1_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 319.170 0.000 319.310 0.350 ;
    END
  END r1_rd_out[8]
  PIN r1_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 330.670 0.000 330.810 0.350 ;
    END
  END r1_rd_out[9]
  PIN r1_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 342.170 0.000 342.310 0.350 ;
    END
  END r1_rd_out[10]
  PIN r1_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 353.670 0.000 353.810 0.350 ;
    END
  END r1_rd_out[11]
  PIN r1_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 365.170 0.000 365.310 0.350 ;
    END
  END r1_rd_out[12]
  PIN r1_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 376.670 0.000 376.810 0.350 ;
    END
  END r1_rd_out[13]
  PIN r1_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 388.170 0.000 388.310 0.350 ;
    END
  END r1_rd_out[14]
  PIN r1_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 399.670 0.000 399.810 0.350 ;
    END
  END r1_rd_out[15]
  PIN r1_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 411.170 0.000 411.310 0.350 ;
    END
  END r1_rd_out[16]
  PIN r1_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 422.670 0.000 422.810 0.350 ;
    END
  END r1_rd_out[17]
  PIN r1_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 434.170 0.000 434.310 0.350 ;
    END
  END r1_rd_out[18]
  PIN r1_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 445.670 0.000 445.810 0.350 ;
    END
  END r1_rd_out[19]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 477.140 6.650 477.940 6.950 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 477.140 12.770 477.940 13.070 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 477.140 18.890 477.940 19.190 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 477.140 25.010 477.940 25.310 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 477.140 31.130 477.940 31.430 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 477.140 37.250 477.940 37.550 ;
    END
  END w0_addr_in[5]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 190.050 4.670 190.400 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 15.110 190.050 15.250 190.400 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 25.690 190.050 25.830 190.400 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 36.270 190.050 36.410 190.400 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 46.850 190.050 46.990 190.400 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 57.430 190.050 57.570 190.400 ;
    END
  END r0_addr_in[5]
  PIN r1_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 58.810 190.050 58.950 190.400 ;
    END
  END r1_addr_in[0]
  PIN r1_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 69.390 190.050 69.530 190.400 ;
    END
  END r1_addr_in[1]
  PIN r1_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 79.970 190.050 80.110 190.400 ;
    END
  END r1_addr_in[2]
  PIN r1_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 90.550 190.050 90.690 190.400 ;
    END
  END r1_addr_in[3]
  PIN r1_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 101.130 190.050 101.270 190.400 ;
    END
  END r1_addr_in[4]
  PIN r1_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 111.710 190.050 111.850 190.400 ;
    END
  END r1_addr_in[5]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 477.140 46.090 477.940 46.390 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 477.140 54.930 477.940 55.230 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 477.140 63.770 477.940 64.070 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 113.090 190.050 113.230 190.400 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 114.470 190.050 114.610 190.400 ;
    END
  END r0_clk
  PIN r1_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 115.850 190.050 115.990 190.400 ;
    END
  END r1_ce_in
  PIN r1_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 117.230 190.050 117.370 190.400 ;
    END
  END r1_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 3.240 6.800 5.960 183.600 ;
      RECT 14.120 6.800 16.840 183.600 ;
      RECT 25.000 6.800 27.720 183.600 ;
      RECT 35.880 6.800 38.600 183.600 ;
      RECT 46.760 6.800 49.480 183.600 ;
      RECT 57.640 6.800 60.360 183.600 ;
      RECT 68.520 6.800 71.240 183.600 ;
      RECT 79.400 6.800 82.120 183.600 ;
      RECT 90.280 6.800 93.000 183.600 ;
      RECT 101.160 6.800 103.880 183.600 ;
      RECT 112.040 6.800 114.760 183.600 ;
      RECT 122.920 6.800 125.640 183.600 ;
      RECT 133.800 6.800 136.520 183.600 ;
      RECT 144.680 6.800 147.400 183.600 ;
      RECT 155.560 6.800 158.280 183.600 ;
      RECT 166.440 6.800 169.160 183.600 ;
      RECT 177.320 6.800 180.040 183.600 ;
      RECT 188.200 6.800 190.920 183.600 ;
      RECT 199.080 6.800 201.800 183.600 ;
      RECT 209.960 6.800 212.680 183.600 ;
      RECT 220.840 6.800 223.560 183.600 ;
      RECT 231.720 6.800 234.440 183.600 ;
      RECT 242.600 6.800 245.320 183.600 ;
      RECT 253.480 6.800 256.200 183.600 ;
      RECT 264.360 6.800 267.080 183.600 ;
      RECT 275.240 6.800 277.960 183.600 ;
      RECT 286.120 6.800 288.840 183.600 ;
      RECT 297.000 6.800 299.720 183.600 ;
      RECT 307.880 6.800 310.600 183.600 ;
      RECT 318.760 6.800 321.480 183.600 ;
      RECT 329.640 6.800 332.360 183.600 ;
      RECT 340.520 6.800 343.240 183.600 ;
      RECT 351.400 6.800 354.120 183.600 ;
      RECT 362.280 6.800 365.000 183.600 ;
      RECT 373.160 6.800 375.880 183.600 ;
      RECT 384.040 6.800 386.760 183.600 ;
      RECT 394.920 6.800 397.640 183.600 ;
      RECT 405.800 6.800 408.520 183.600 ;
      RECT 416.680 6.800 419.400 183.600 ;
      RECT 427.560 6.800 430.280 183.600 ;
      RECT 438.440 6.800 441.160 183.600 ;
      RECT 449.320 6.800 452.040 183.600 ;
      RECT 460.200 6.800 462.920 183.600 ;
      RECT 471.080 6.800 473.800 183.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 8.680 6.800 11.400 183.600 ;
      RECT 19.560 6.800 22.280 183.600 ;
      RECT 30.440 6.800 33.160 183.600 ;
      RECT 41.320 6.800 44.040 183.600 ;
      RECT 52.200 6.800 54.920 183.600 ;
      RECT 63.080 6.800 65.800 183.600 ;
      RECT 73.960 6.800 76.680 183.600 ;
      RECT 84.840 6.800 87.560 183.600 ;
      RECT 95.720 6.800 98.440 183.600 ;
      RECT 106.600 6.800 109.320 183.600 ;
      RECT 117.480 6.800 120.200 183.600 ;
      RECT 128.360 6.800 131.080 183.600 ;
      RECT 139.240 6.800 141.960 183.600 ;
      RECT 150.120 6.800 152.840 183.600 ;
      RECT 161.000 6.800 163.720 183.600 ;
      RECT 171.880 6.800 174.600 183.600 ;
      RECT 182.760 6.800 185.480 183.600 ;
      RECT 193.640 6.800 196.360 183.600 ;
      RECT 204.520 6.800 207.240 183.600 ;
      RECT 215.400 6.800 218.120 183.600 ;
      RECT 226.280 6.800 229.000 183.600 ;
      RECT 237.160 6.800 239.880 183.600 ;
      RECT 248.040 6.800 250.760 183.600 ;
      RECT 258.920 6.800 261.640 183.600 ;
      RECT 269.800 6.800 272.520 183.600 ;
      RECT 280.680 6.800 283.400 183.600 ;
      RECT 291.560 6.800 294.280 183.600 ;
      RECT 302.440 6.800 305.160 183.600 ;
      RECT 313.320 6.800 316.040 183.600 ;
      RECT 324.200 6.800 326.920 183.600 ;
      RECT 335.080 6.800 337.800 183.600 ;
      RECT 345.960 6.800 348.680 183.600 ;
      RECT 356.840 6.800 359.560 183.600 ;
      RECT 367.720 6.800 370.440 183.600 ;
      RECT 378.600 6.800 381.320 183.600 ;
      RECT 389.480 6.800 392.200 183.600 ;
      RECT 400.360 6.800 403.080 183.600 ;
      RECT 411.240 6.800 413.960 183.600 ;
      RECT 422.120 6.800 424.840 183.600 ;
      RECT 433.000 6.800 435.720 183.600 ;
      RECT 443.880 6.800 446.600 183.600 ;
      RECT 454.760 6.800 457.480 183.600 ;
      RECT 465.640 6.800 468.360 183.600 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 477.940 190.400 ;
    LAYER met2 ;
    RECT 0 0 477.940 190.400 ;
    LAYER met3 ;
    RECT 0.800 0 477.940 190.400 ;
    LAYER met4 ;
    RECT 0 0 477.940 6.800 ;
    RECT 0 183.600 477.940 190.400 ;
    RECT 0.000 6.800 3.240 183.600 ;
    RECT 5.960 6.800 8.680 183.600 ;
    RECT 11.400 6.800 14.120 183.600 ;
    RECT 16.840 6.800 19.560 183.600 ;
    RECT 22.280 6.800 25.000 183.600 ;
    RECT 27.720 6.800 30.440 183.600 ;
    RECT 33.160 6.800 35.880 183.600 ;
    RECT 38.600 6.800 41.320 183.600 ;
    RECT 44.040 6.800 46.760 183.600 ;
    RECT 49.480 6.800 52.200 183.600 ;
    RECT 54.920 6.800 57.640 183.600 ;
    RECT 60.360 6.800 63.080 183.600 ;
    RECT 65.800 6.800 68.520 183.600 ;
    RECT 71.240 6.800 73.960 183.600 ;
    RECT 76.680 6.800 79.400 183.600 ;
    RECT 82.120 6.800 84.840 183.600 ;
    RECT 87.560 6.800 90.280 183.600 ;
    RECT 93.000 6.800 95.720 183.600 ;
    RECT 98.440 6.800 101.160 183.600 ;
    RECT 103.880 6.800 106.600 183.600 ;
    RECT 109.320 6.800 112.040 183.600 ;
    RECT 114.760 6.800 117.480 183.600 ;
    RECT 120.200 6.800 122.920 183.600 ;
    RECT 125.640 6.800 128.360 183.600 ;
    RECT 131.080 6.800 133.800 183.600 ;
    RECT 136.520 6.800 139.240 183.600 ;
    RECT 141.960 6.800 144.680 183.600 ;
    RECT 147.400 6.800 150.120 183.600 ;
    RECT 152.840 6.800 155.560 183.600 ;
    RECT 158.280 6.800 161.000 183.600 ;
    RECT 163.720 6.800 166.440 183.600 ;
    RECT 169.160 6.800 171.880 183.600 ;
    RECT 174.600 6.800 177.320 183.600 ;
    RECT 180.040 6.800 182.760 183.600 ;
    RECT 185.480 6.800 188.200 183.600 ;
    RECT 190.920 6.800 193.640 183.600 ;
    RECT 196.360 6.800 199.080 183.600 ;
    RECT 201.800 6.800 204.520 183.600 ;
    RECT 207.240 6.800 209.960 183.600 ;
    RECT 212.680 6.800 215.400 183.600 ;
    RECT 218.120 6.800 220.840 183.600 ;
    RECT 223.560 6.800 226.280 183.600 ;
    RECT 229.000 6.800 231.720 183.600 ;
    RECT 234.440 6.800 237.160 183.600 ;
    RECT 239.880 6.800 242.600 183.600 ;
    RECT 245.320 6.800 248.040 183.600 ;
    RECT 250.760 6.800 253.480 183.600 ;
    RECT 256.200 6.800 258.920 183.600 ;
    RECT 261.640 6.800 264.360 183.600 ;
    RECT 267.080 6.800 269.800 183.600 ;
    RECT 272.520 6.800 275.240 183.600 ;
    RECT 277.960 6.800 280.680 183.600 ;
    RECT 283.400 6.800 286.120 183.600 ;
    RECT 288.840 6.800 291.560 183.600 ;
    RECT 294.280 6.800 297.000 183.600 ;
    RECT 299.720 6.800 302.440 183.600 ;
    RECT 305.160 6.800 307.880 183.600 ;
    RECT 310.600 6.800 313.320 183.600 ;
    RECT 316.040 6.800 318.760 183.600 ;
    RECT 321.480 6.800 324.200 183.600 ;
    RECT 326.920 6.800 329.640 183.600 ;
    RECT 332.360 6.800 335.080 183.600 ;
    RECT 337.800 6.800 340.520 183.600 ;
    RECT 343.240 6.800 345.960 183.600 ;
    RECT 348.680 6.800 351.400 183.600 ;
    RECT 354.120 6.800 356.840 183.600 ;
    RECT 359.560 6.800 362.280 183.600 ;
    RECT 365.000 6.800 367.720 183.600 ;
    RECT 370.440 6.800 373.160 183.600 ;
    RECT 375.880 6.800 378.600 183.600 ;
    RECT 381.320 6.800 384.040 183.600 ;
    RECT 386.760 6.800 389.480 183.600 ;
    RECT 392.200 6.800 394.920 183.600 ;
    RECT 397.640 6.800 400.360 183.600 ;
    RECT 403.080 6.800 405.800 183.600 ;
    RECT 408.520 6.800 411.240 183.600 ;
    RECT 413.960 6.800 416.680 183.600 ;
    RECT 419.400 6.800 422.120 183.600 ;
    RECT 424.840 6.800 427.560 183.600 ;
    RECT 430.280 6.800 433.000 183.600 ;
    RECT 435.720 6.800 438.440 183.600 ;
    RECT 441.160 6.800 443.880 183.600 ;
    RECT 446.600 6.800 449.320 183.600 ;
    RECT 452.040 6.800 454.760 183.600 ;
    RECT 457.480 6.800 460.200 183.600 ;
    RECT 462.920 6.800 465.640 183.600 ;
    RECT 468.360 6.800 471.080 183.600 ;
    RECT 473.800 6.800 477.940 183.600 ;
    LAYER OVERLAP ;
    RECT 0 0 477.940 190.400 ;
  END
END fakeram_20x64_2r1w

END LIBRARY
