VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_20x64_1r1w
  FOREIGN fakeram_20x64_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 376.280 BY 138.720 ;
  CLASS BLOCK ;
  PIN w0_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 6.650 0.800 6.950 ;
    END
  END w0_mask_in[0]
  PIN w0_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 9.370 0.800 9.670 ;
    END
  END w0_mask_in[1]
  PIN w0_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 12.090 0.800 12.390 ;
    END
  END w0_mask_in[2]
  PIN w0_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.810 0.800 15.110 ;
    END
  END w0_mask_in[3]
  PIN w0_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 17.530 0.800 17.830 ;
    END
  END w0_mask_in[4]
  PIN w0_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.250 0.800 20.550 ;
    END
  END w0_mask_in[5]
  PIN w0_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.970 0.800 23.270 ;
    END
  END w0_mask_in[6]
  PIN w0_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 25.690 0.800 25.990 ;
    END
  END w0_mask_in[7]
  PIN w0_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 28.410 0.800 28.710 ;
    END
  END w0_mask_in[8]
  PIN w0_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.130 0.800 31.430 ;
    END
  END w0_mask_in[9]
  PIN w0_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 33.850 0.800 34.150 ;
    END
  END w0_mask_in[10]
  PIN w0_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 36.570 0.800 36.870 ;
    END
  END w0_mask_in[11]
  PIN w0_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.290 0.800 39.590 ;
    END
  END w0_mask_in[12]
  PIN w0_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 42.010 0.800 42.310 ;
    END
  END w0_mask_in[13]
  PIN w0_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 44.730 0.800 45.030 ;
    END
  END w0_mask_in[14]
  PIN w0_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 47.450 0.800 47.750 ;
    END
  END w0_mask_in[15]
  PIN w0_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 50.170 0.800 50.470 ;
    END
  END w0_mask_in[16]
  PIN w0_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 52.890 0.800 53.190 ;
    END
  END w0_mask_in[17]
  PIN w0_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.610 0.800 55.910 ;
    END
  END w0_mask_in[18]
  PIN w0_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 58.330 0.800 58.630 ;
    END
  END w0_mask_in[19]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 66.490 0.800 66.790 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 69.210 0.800 69.510 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.930 0.800 72.230 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 74.650 0.800 74.950 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 77.370 0.800 77.670 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 80.090 0.800 80.390 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 82.810 0.800 83.110 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 85.530 0.800 85.830 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 88.250 0.800 88.550 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 90.970 0.800 91.270 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 93.690 0.800 93.990 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 96.410 0.800 96.710 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 99.130 0.800 99.430 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 101.850 0.800 102.150 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 104.570 0.800 104.870 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 107.290 0.800 107.590 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 110.010 0.800 110.310 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 112.730 0.800 113.030 ;
    END
  END w0_wd_in[17]
  PIN w0_wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 115.450 0.800 115.750 ;
    END
  END w0_wd_in[18]
  PIN w0_wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 118.170 0.800 118.470 ;
    END
  END w0_wd_in[19]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 0.000 4.670 0.350 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 22.470 0.000 22.610 0.350 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 40.410 0.000 40.550 0.350 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 58.350 0.000 58.490 0.350 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 76.290 0.000 76.430 0.350 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 94.230 0.000 94.370 0.350 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 112.170 0.000 112.310 0.350 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 130.110 0.000 130.250 0.350 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 148.050 0.000 148.190 0.350 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 165.990 0.000 166.130 0.350 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 183.930 0.000 184.070 0.350 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 201.870 0.000 202.010 0.350 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 219.810 0.000 219.950 0.350 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 237.750 0.000 237.890 0.350 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 255.690 0.000 255.830 0.350 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 273.630 0.000 273.770 0.350 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 291.570 0.000 291.710 0.350 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 309.510 0.000 309.650 0.350 ;
    END
  END r0_rd_out[17]
  PIN r0_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 327.450 0.000 327.590 0.350 ;
    END
  END r0_rd_out[18]
  PIN r0_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 345.390 0.000 345.530 0.350 ;
    END
  END r0_rd_out[19]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 6.650 376.280 6.950 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 11.410 376.280 11.710 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 16.170 376.280 16.470 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 20.930 376.280 21.230 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 25.690 376.280 25.990 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 30.450 376.280 30.750 ;
    END
  END w0_addr_in[5]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 138.370 4.670 138.720 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 21.090 138.370 21.230 138.720 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 37.650 138.370 37.790 138.720 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 54.210 138.370 54.350 138.720 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 70.770 138.370 70.910 138.720 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 87.330 138.370 87.470 138.720 ;
    END
  END r0_addr_in[5]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 37.930 376.280 38.230 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 45.410 376.280 45.710 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 375.480 52.890 376.280 53.190 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 88.250 138.370 88.390 138.720 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 89.170 138.370 89.310 138.720 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 3.240 6.800 5.960 131.920 ;
      RECT 14.120 6.800 16.840 131.920 ;
      RECT 25.000 6.800 27.720 131.920 ;
      RECT 35.880 6.800 38.600 131.920 ;
      RECT 46.760 6.800 49.480 131.920 ;
      RECT 57.640 6.800 60.360 131.920 ;
      RECT 68.520 6.800 71.240 131.920 ;
      RECT 79.400 6.800 82.120 131.920 ;
      RECT 90.280 6.800 93.000 131.920 ;
      RECT 101.160 6.800 103.880 131.920 ;
      RECT 112.040 6.800 114.760 131.920 ;
      RECT 122.920 6.800 125.640 131.920 ;
      RECT 133.800 6.800 136.520 131.920 ;
      RECT 144.680 6.800 147.400 131.920 ;
      RECT 155.560 6.800 158.280 131.920 ;
      RECT 166.440 6.800 169.160 131.920 ;
      RECT 177.320 6.800 180.040 131.920 ;
      RECT 188.200 6.800 190.920 131.920 ;
      RECT 199.080 6.800 201.800 131.920 ;
      RECT 209.960 6.800 212.680 131.920 ;
      RECT 220.840 6.800 223.560 131.920 ;
      RECT 231.720 6.800 234.440 131.920 ;
      RECT 242.600 6.800 245.320 131.920 ;
      RECT 253.480 6.800 256.200 131.920 ;
      RECT 264.360 6.800 267.080 131.920 ;
      RECT 275.240 6.800 277.960 131.920 ;
      RECT 286.120 6.800 288.840 131.920 ;
      RECT 297.000 6.800 299.720 131.920 ;
      RECT 307.880 6.800 310.600 131.920 ;
      RECT 318.760 6.800 321.480 131.920 ;
      RECT 329.640 6.800 332.360 131.920 ;
      RECT 340.520 6.800 343.240 131.920 ;
      RECT 351.400 6.800 354.120 131.920 ;
      RECT 362.280 6.800 365.000 131.920 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 8.680 6.800 11.400 131.920 ;
      RECT 19.560 6.800 22.280 131.920 ;
      RECT 30.440 6.800 33.160 131.920 ;
      RECT 41.320 6.800 44.040 131.920 ;
      RECT 52.200 6.800 54.920 131.920 ;
      RECT 63.080 6.800 65.800 131.920 ;
      RECT 73.960 6.800 76.680 131.920 ;
      RECT 84.840 6.800 87.560 131.920 ;
      RECT 95.720 6.800 98.440 131.920 ;
      RECT 106.600 6.800 109.320 131.920 ;
      RECT 117.480 6.800 120.200 131.920 ;
      RECT 128.360 6.800 131.080 131.920 ;
      RECT 139.240 6.800 141.960 131.920 ;
      RECT 150.120 6.800 152.840 131.920 ;
      RECT 161.000 6.800 163.720 131.920 ;
      RECT 171.880 6.800 174.600 131.920 ;
      RECT 182.760 6.800 185.480 131.920 ;
      RECT 193.640 6.800 196.360 131.920 ;
      RECT 204.520 6.800 207.240 131.920 ;
      RECT 215.400 6.800 218.120 131.920 ;
      RECT 226.280 6.800 229.000 131.920 ;
      RECT 237.160 6.800 239.880 131.920 ;
      RECT 248.040 6.800 250.760 131.920 ;
      RECT 258.920 6.800 261.640 131.920 ;
      RECT 269.800 6.800 272.520 131.920 ;
      RECT 280.680 6.800 283.400 131.920 ;
      RECT 291.560 6.800 294.280 131.920 ;
      RECT 302.440 6.800 305.160 131.920 ;
      RECT 313.320 6.800 316.040 131.920 ;
      RECT 324.200 6.800 326.920 131.920 ;
      RECT 335.080 6.800 337.800 131.920 ;
      RECT 345.960 6.800 348.680 131.920 ;
      RECT 356.840 6.800 359.560 131.920 ;
      RECT 367.720 6.800 370.440 131.920 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 376.280 138.720 ;
    LAYER met2 ;
    RECT 0 0 376.280 138.720 ;
    LAYER met3 ;
    RECT 0.800 0 376.280 138.720 ;
    LAYER met4 ;
    RECT 0 0 376.280 6.800 ;
    RECT 0 131.920 376.280 138.720 ;
    RECT 0.000 6.800 3.240 131.920 ;
    RECT 5.960 6.800 8.680 131.920 ;
    RECT 11.400 6.800 14.120 131.920 ;
    RECT 16.840 6.800 19.560 131.920 ;
    RECT 22.280 6.800 25.000 131.920 ;
    RECT 27.720 6.800 30.440 131.920 ;
    RECT 33.160 6.800 35.880 131.920 ;
    RECT 38.600 6.800 41.320 131.920 ;
    RECT 44.040 6.800 46.760 131.920 ;
    RECT 49.480 6.800 52.200 131.920 ;
    RECT 54.920 6.800 57.640 131.920 ;
    RECT 60.360 6.800 63.080 131.920 ;
    RECT 65.800 6.800 68.520 131.920 ;
    RECT 71.240 6.800 73.960 131.920 ;
    RECT 76.680 6.800 79.400 131.920 ;
    RECT 82.120 6.800 84.840 131.920 ;
    RECT 87.560 6.800 90.280 131.920 ;
    RECT 93.000 6.800 95.720 131.920 ;
    RECT 98.440 6.800 101.160 131.920 ;
    RECT 103.880 6.800 106.600 131.920 ;
    RECT 109.320 6.800 112.040 131.920 ;
    RECT 114.760 6.800 117.480 131.920 ;
    RECT 120.200 6.800 122.920 131.920 ;
    RECT 125.640 6.800 128.360 131.920 ;
    RECT 131.080 6.800 133.800 131.920 ;
    RECT 136.520 6.800 139.240 131.920 ;
    RECT 141.960 6.800 144.680 131.920 ;
    RECT 147.400 6.800 150.120 131.920 ;
    RECT 152.840 6.800 155.560 131.920 ;
    RECT 158.280 6.800 161.000 131.920 ;
    RECT 163.720 6.800 166.440 131.920 ;
    RECT 169.160 6.800 171.880 131.920 ;
    RECT 174.600 6.800 177.320 131.920 ;
    RECT 180.040 6.800 182.760 131.920 ;
    RECT 185.480 6.800 188.200 131.920 ;
    RECT 190.920 6.800 193.640 131.920 ;
    RECT 196.360 6.800 199.080 131.920 ;
    RECT 201.800 6.800 204.520 131.920 ;
    RECT 207.240 6.800 209.960 131.920 ;
    RECT 212.680 6.800 215.400 131.920 ;
    RECT 218.120 6.800 220.840 131.920 ;
    RECT 223.560 6.800 226.280 131.920 ;
    RECT 229.000 6.800 231.720 131.920 ;
    RECT 234.440 6.800 237.160 131.920 ;
    RECT 239.880 6.800 242.600 131.920 ;
    RECT 245.320 6.800 248.040 131.920 ;
    RECT 250.760 6.800 253.480 131.920 ;
    RECT 256.200 6.800 258.920 131.920 ;
    RECT 261.640 6.800 264.360 131.920 ;
    RECT 267.080 6.800 269.800 131.920 ;
    RECT 272.520 6.800 275.240 131.920 ;
    RECT 277.960 6.800 280.680 131.920 ;
    RECT 283.400 6.800 286.120 131.920 ;
    RECT 288.840 6.800 291.560 131.920 ;
    RECT 294.280 6.800 297.000 131.920 ;
    RECT 299.720 6.800 302.440 131.920 ;
    RECT 305.160 6.800 307.880 131.920 ;
    RECT 310.600 6.800 313.320 131.920 ;
    RECT 316.040 6.800 318.760 131.920 ;
    RECT 321.480 6.800 324.200 131.920 ;
    RECT 326.920 6.800 329.640 131.920 ;
    RECT 332.360 6.800 335.080 131.920 ;
    RECT 337.800 6.800 340.520 131.920 ;
    RECT 343.240 6.800 345.960 131.920 ;
    RECT 348.680 6.800 351.400 131.920 ;
    RECT 354.120 6.800 356.840 131.920 ;
    RECT 359.560 6.800 362.280 131.920 ;
    RECT 365.000 6.800 367.720 131.920 ;
    RECT 370.440 6.800 376.280 131.920 ;
    LAYER OVERLAP ;
    RECT 0 0 376.280 138.720 ;
  END
END fakeram_20x64_1r1w

END LIBRARY
