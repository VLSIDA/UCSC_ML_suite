VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO liteeth_1rw1r_32w384d_8_sram
  FOREIGN liteeth_1rw1r_32w384d_8_sram 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 114.000 BY 256.200 ;
  CLASS BLOCK ;
  PIN w_mask_rw1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 -0.595 0.070 -0.525 ;
    END
  END w_mask_rw1[0]
  PIN w_mask_rw1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.505 0.070 1.575 ;
    END
  END w_mask_rw1[1]
  PIN w_mask_rw1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.605 0.070 3.675 ;
    END
  END w_mask_rw1[2]
  PIN w_mask_rw1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.705 0.070 5.775 ;
    END
  END w_mask_rw1[3]
  PIN w_mask_rw1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.805 0.070 7.875 ;
    END
  END w_mask_rw1[4]
  PIN w_mask_rw1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.905 0.070 9.975 ;
    END
  END w_mask_rw1[5]
  PIN w_mask_rw1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.005 0.070 12.075 ;
    END
  END w_mask_rw1[6]
  PIN w_mask_rw1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.105 0.070 14.175 ;
    END
  END w_mask_rw1[7]
  PIN w_mask_rw1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.205 0.070 16.275 ;
    END
  END w_mask_rw1[8]
  PIN w_mask_rw1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.305 0.070 18.375 ;
    END
  END w_mask_rw1[9]
  PIN w_mask_rw1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.405 0.070 20.475 ;
    END
  END w_mask_rw1[10]
  PIN w_mask_rw1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.505 0.070 22.575 ;
    END
  END w_mask_rw1[11]
  PIN w_mask_rw1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.605 0.070 24.675 ;
    END
  END w_mask_rw1[12]
  PIN w_mask_rw1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.705 0.070 26.775 ;
    END
  END w_mask_rw1[13]
  PIN w_mask_rw1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.805 0.070 28.875 ;
    END
  END w_mask_rw1[14]
  PIN w_mask_rw1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.905 0.070 30.975 ;
    END
  END w_mask_rw1[15]
  PIN w_mask_rw1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.005 0.070 33.075 ;
    END
  END w_mask_rw1[16]
  PIN w_mask_rw1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.105 0.070 35.175 ;
    END
  END w_mask_rw1[17]
  PIN w_mask_rw1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.205 0.070 37.275 ;
    END
  END w_mask_rw1[18]
  PIN w_mask_rw1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.305 0.070 39.375 ;
    END
  END w_mask_rw1[19]
  PIN w_mask_rw1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.405 0.070 41.475 ;
    END
  END w_mask_rw1[20]
  PIN w_mask_rw1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.505 0.070 43.575 ;
    END
  END w_mask_rw1[21]
  PIN w_mask_rw1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.605 0.070 45.675 ;
    END
  END w_mask_rw1[22]
  PIN w_mask_rw1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.705 0.070 47.775 ;
    END
  END w_mask_rw1[23]
  PIN w_mask_rw1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.805 0.070 49.875 ;
    END
  END w_mask_rw1[24]
  PIN w_mask_rw1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.905 0.070 51.975 ;
    END
  END w_mask_rw1[25]
  PIN w_mask_rw1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.005 0.070 54.075 ;
    END
  END w_mask_rw1[26]
  PIN w_mask_rw1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.105 0.070 56.175 ;
    END
  END w_mask_rw1[27]
  PIN w_mask_rw1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.205 0.070 58.275 ;
    END
  END w_mask_rw1[28]
  PIN w_mask_rw1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.305 0.070 60.375 ;
    END
  END w_mask_rw1[29]
  PIN w_mask_rw1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.405 0.070 62.475 ;
    END
  END w_mask_rw1[30]
  PIN w_mask_rw1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.505 0.070 64.575 ;
    END
  END w_mask_rw1[31]
  PIN rd_out_rw1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.645 0.070 64.715 ;
    END
  END rd_out_rw1[0]
  PIN rd_out_rw1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.745 0.070 66.815 ;
    END
  END rd_out_rw1[1]
  PIN rd_out_rw1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END rd_out_rw1[2]
  PIN rd_out_rw1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END rd_out_rw1[3]
  PIN rd_out_rw1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END rd_out_rw1[4]
  PIN rd_out_rw1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END rd_out_rw1[5]
  PIN rd_out_rw1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END rd_out_rw1[6]
  PIN rd_out_rw1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END rd_out_rw1[7]
  PIN rd_out_rw1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END rd_out_rw1[8]
  PIN rd_out_rw1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END rd_out_rw1[9]
  PIN rd_out_rw1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END rd_out_rw1[10]
  PIN rd_out_rw1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.745 0.070 87.815 ;
    END
  END rd_out_rw1[11]
  PIN rd_out_rw1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.845 0.070 89.915 ;
    END
  END rd_out_rw1[12]
  PIN rd_out_rw1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.945 0.070 92.015 ;
    END
  END rd_out_rw1[13]
  PIN rd_out_rw1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.045 0.070 94.115 ;
    END
  END rd_out_rw1[14]
  PIN rd_out_rw1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.145 0.070 96.215 ;
    END
  END rd_out_rw1[15]
  PIN rd_out_rw1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.245 0.070 98.315 ;
    END
  END rd_out_rw1[16]
  PIN rd_out_rw1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.345 0.070 100.415 ;
    END
  END rd_out_rw1[17]
  PIN rd_out_rw1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.445 0.070 102.515 ;
    END
  END rd_out_rw1[18]
  PIN rd_out_rw1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.545 0.070 104.615 ;
    END
  END rd_out_rw1[19]
  PIN rd_out_rw1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.645 0.070 106.715 ;
    END
  END rd_out_rw1[20]
  PIN rd_out_rw1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.745 0.070 108.815 ;
    END
  END rd_out_rw1[21]
  PIN rd_out_rw1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.845 0.070 110.915 ;
    END
  END rd_out_rw1[22]
  PIN rd_out_rw1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.945 0.070 113.015 ;
    END
  END rd_out_rw1[23]
  PIN rd_out_rw1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.045 0.070 115.115 ;
    END
  END rd_out_rw1[24]
  PIN rd_out_rw1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.145 0.070 117.215 ;
    END
  END rd_out_rw1[25]
  PIN rd_out_rw1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.245 0.070 119.315 ;
    END
  END rd_out_rw1[26]
  PIN rd_out_rw1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.345 0.070 121.415 ;
    END
  END rd_out_rw1[27]
  PIN rd_out_rw1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.445 0.070 123.515 ;
    END
  END rd_out_rw1[28]
  PIN rd_out_rw1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.545 0.070 125.615 ;
    END
  END rd_out_rw1[29]
  PIN rd_out_rw1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.645 0.070 127.715 ;
    END
  END rd_out_rw1[30]
  PIN rd_out_rw1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.745 0.070 129.815 ;
    END
  END rd_out_rw1[31]
  PIN rd_out_r1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.885 0.070 129.955 ;
    END
  END rd_out_r1[0]
  PIN rd_out_r1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.985 0.070 132.055 ;
    END
  END rd_out_r1[1]
  PIN rd_out_r1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.085 0.070 134.155 ;
    END
  END rd_out_r1[2]
  PIN rd_out_r1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.185 0.070 136.255 ;
    END
  END rd_out_r1[3]
  PIN rd_out_r1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.285 0.070 138.355 ;
    END
  END rd_out_r1[4]
  PIN rd_out_r1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.385 0.070 140.455 ;
    END
  END rd_out_r1[5]
  PIN rd_out_r1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.485 0.070 142.555 ;
    END
  END rd_out_r1[6]
  PIN rd_out_r1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.585 0.070 144.655 ;
    END
  END rd_out_r1[7]
  PIN rd_out_r1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.685 0.070 146.755 ;
    END
  END rd_out_r1[8]
  PIN rd_out_r1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.785 0.070 148.855 ;
    END
  END rd_out_r1[9]
  PIN rd_out_r1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.885 0.070 150.955 ;
    END
  END rd_out_r1[10]
  PIN rd_out_r1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.985 0.070 153.055 ;
    END
  END rd_out_r1[11]
  PIN rd_out_r1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.085 0.070 155.155 ;
    END
  END rd_out_r1[12]
  PIN rd_out_r1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.185 0.070 157.255 ;
    END
  END rd_out_r1[13]
  PIN rd_out_r1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.285 0.070 159.355 ;
    END
  END rd_out_r1[14]
  PIN rd_out_r1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.385 0.070 161.455 ;
    END
  END rd_out_r1[15]
  PIN rd_out_r1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.485 0.070 163.555 ;
    END
  END rd_out_r1[16]
  PIN rd_out_r1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.585 0.070 165.655 ;
    END
  END rd_out_r1[17]
  PIN rd_out_r1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.685 0.070 167.755 ;
    END
  END rd_out_r1[18]
  PIN rd_out_r1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.785 0.070 169.855 ;
    END
  END rd_out_r1[19]
  PIN rd_out_r1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.885 0.070 171.955 ;
    END
  END rd_out_r1[20]
  PIN rd_out_r1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.985 0.070 174.055 ;
    END
  END rd_out_r1[21]
  PIN rd_out_r1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.085 0.070 176.155 ;
    END
  END rd_out_r1[22]
  PIN rd_out_r1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.185 0.070 178.255 ;
    END
  END rd_out_r1[23]
  PIN rd_out_r1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.285 0.070 180.355 ;
    END
  END rd_out_r1[24]
  PIN rd_out_r1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.385 0.070 182.455 ;
    END
  END rd_out_r1[25]
  PIN rd_out_r1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.485 0.070 184.555 ;
    END
  END rd_out_r1[26]
  PIN rd_out_r1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.585 0.070 186.655 ;
    END
  END rd_out_r1[27]
  PIN rd_out_r1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.685 0.070 188.755 ;
    END
  END rd_out_r1[28]
  PIN rd_out_r1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.785 0.070 190.855 ;
    END
  END rd_out_r1[29]
  PIN rd_out_r1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.885 0.070 192.955 ;
    END
  END rd_out_r1[30]
  PIN rd_out_r1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.985 0.070 195.055 ;
    END
  END rd_out_r1[31]
  PIN wd_in_rw1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.125 0.070 195.195 ;
    END
  END wd_in_rw1[0]
  PIN wd_in_rw1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.225 0.070 197.295 ;
    END
  END wd_in_rw1[1]
  PIN wd_in_rw1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.325 0.070 199.395 ;
    END
  END wd_in_rw1[2]
  PIN wd_in_rw1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.425 0.070 201.495 ;
    END
  END wd_in_rw1[3]
  PIN wd_in_rw1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.525 0.070 203.595 ;
    END
  END wd_in_rw1[4]
  PIN wd_in_rw1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.625 0.070 205.695 ;
    END
  END wd_in_rw1[5]
  PIN wd_in_rw1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.725 0.070 207.795 ;
    END
  END wd_in_rw1[6]
  PIN wd_in_rw1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.825 0.070 209.895 ;
    END
  END wd_in_rw1[7]
  PIN wd_in_rw1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.925 0.070 211.995 ;
    END
  END wd_in_rw1[8]
  PIN wd_in_rw1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.025 0.070 214.095 ;
    END
  END wd_in_rw1[9]
  PIN wd_in_rw1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.125 0.070 216.195 ;
    END
  END wd_in_rw1[10]
  PIN wd_in_rw1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.225 0.070 218.295 ;
    END
  END wd_in_rw1[11]
  PIN wd_in_rw1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.325 0.070 220.395 ;
    END
  END wd_in_rw1[12]
  PIN wd_in_rw1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.425 0.070 222.495 ;
    END
  END wd_in_rw1[13]
  PIN wd_in_rw1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.525 0.070 224.595 ;
    END
  END wd_in_rw1[14]
  PIN wd_in_rw1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.625 0.070 226.695 ;
    END
  END wd_in_rw1[15]
  PIN wd_in_rw1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.725 0.070 228.795 ;
    END
  END wd_in_rw1[16]
  PIN wd_in_rw1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.825 0.070 230.895 ;
    END
  END wd_in_rw1[17]
  PIN wd_in_rw1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.925 0.070 232.995 ;
    END
  END wd_in_rw1[18]
  PIN wd_in_rw1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.025 0.070 235.095 ;
    END
  END wd_in_rw1[19]
  PIN wd_in_rw1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.125 0.070 237.195 ;
    END
  END wd_in_rw1[20]
  PIN wd_in_rw1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.225 0.070 239.295 ;
    END
  END wd_in_rw1[21]
  PIN wd_in_rw1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.325 0.070 241.395 ;
    END
  END wd_in_rw1[22]
  PIN wd_in_rw1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.425 0.070 243.495 ;
    END
  END wd_in_rw1[23]
  PIN wd_in_rw1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 245.525 0.070 245.595 ;
    END
  END wd_in_rw1[24]
  PIN wd_in_rw1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.625 0.070 247.695 ;
    END
  END wd_in_rw1[25]
  PIN wd_in_rw1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.725 0.070 249.795 ;
    END
  END wd_in_rw1[26]
  PIN wd_in_rw1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.825 0.070 251.895 ;
    END
  END wd_in_rw1[27]
  PIN wd_in_rw1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.925 0.070 253.995 ;
    END
  END wd_in_rw1[28]
  PIN wd_in_rw1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.025 0.070 256.095 ;
    END
  END wd_in_rw1[29]
  PIN wd_in_rw1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.125 0.070 258.195 ;
    END
  END wd_in_rw1[30]
  PIN wd_in_rw1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.225 0.070 260.295 ;
    END
  END wd_in_rw1[31]
  PIN addr_rw1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.365 0.070 260.435 ;
    END
  END addr_rw1[0]
  PIN addr_rw1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.465 0.070 262.535 ;
    END
  END addr_rw1[1]
  PIN addr_rw1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.565 0.070 264.635 ;
    END
  END addr_rw1[2]
  PIN addr_rw1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.665 0.070 266.735 ;
    END
  END addr_rw1[3]
  PIN addr_rw1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.765 0.070 268.835 ;
    END
  END addr_rw1[4]
  PIN addr_rw1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.865 0.070 270.935 ;
    END
  END addr_rw1[5]
  PIN addr_rw1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.965 0.070 273.035 ;
    END
  END addr_rw1[6]
  PIN addr_rw1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.065 0.070 275.135 ;
    END
  END addr_rw1[7]
  PIN addr_rw1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.165 0.070 277.235 ;
    END
  END addr_rw1[8]
  PIN addr_r1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.305 0.070 277.375 ;
    END
  END addr_r1[0]
  PIN addr_r1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.405 0.070 279.475 ;
    END
  END addr_r1[1]
  PIN addr_r1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.505 0.070 281.575 ;
    END
  END addr_r1[2]
  PIN addr_r1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.605 0.070 283.675 ;
    END
  END addr_r1[3]
  PIN addr_r1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.705 0.070 285.775 ;
    END
  END addr_r1[4]
  PIN addr_r1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.805 0.070 287.875 ;
    END
  END addr_r1[5]
  PIN addr_r1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.905 0.070 289.975 ;
    END
  END addr_r1[6]
  PIN addr_r1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.005 0.070 292.075 ;
    END
  END addr_r1[7]
  PIN addr_r1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.105 0.070 294.175 ;
    END
  END addr_r1[8]
  PIN we_in_rw1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.245 0.070 294.315 ;
    END
  END we_in_rw1
  PIN ce_rw1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.425 0.070 292.495 ;
    END
  END ce_rw1
  PIN ce_r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.605 0.070 290.675 ;
    END
  END ce_r1
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.745 0.070 290.815 ;
    END
  END clk0
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.845 0.070 292.915 ;
    END
  END clk1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 254.800 ;
      RECT 3.500 1.400 3.780 254.800 ;
      RECT 5.740 1.400 6.020 254.800 ;
      RECT 7.980 1.400 8.260 254.800 ;
      RECT 10.220 1.400 10.500 254.800 ;
      RECT 12.460 1.400 12.740 254.800 ;
      RECT 14.700 1.400 14.980 254.800 ;
      RECT 16.940 1.400 17.220 254.800 ;
      RECT 19.180 1.400 19.460 254.800 ;
      RECT 21.420 1.400 21.700 254.800 ;
      RECT 23.660 1.400 23.940 254.800 ;
      RECT 25.900 1.400 26.180 254.800 ;
      RECT 28.140 1.400 28.420 254.800 ;
      RECT 30.380 1.400 30.660 254.800 ;
      RECT 32.620 1.400 32.900 254.800 ;
      RECT 34.860 1.400 35.140 254.800 ;
      RECT 37.100 1.400 37.380 254.800 ;
      RECT 39.340 1.400 39.620 254.800 ;
      RECT 41.580 1.400 41.860 254.800 ;
      RECT 43.820 1.400 44.100 254.800 ;
      RECT 46.060 1.400 46.340 254.800 ;
      RECT 48.300 1.400 48.580 254.800 ;
      RECT 50.540 1.400 50.820 254.800 ;
      RECT 52.780 1.400 53.060 254.800 ;
      RECT 55.020 1.400 55.300 254.800 ;
      RECT 57.260 1.400 57.540 254.800 ;
      RECT 59.500 1.400 59.780 254.800 ;
      RECT 61.740 1.400 62.020 254.800 ;
      RECT 63.980 1.400 64.260 254.800 ;
      RECT 66.220 1.400 66.500 254.800 ;
      RECT 68.460 1.400 68.740 254.800 ;
      RECT 70.700 1.400 70.980 254.800 ;
      RECT 72.940 1.400 73.220 254.800 ;
      RECT 75.180 1.400 75.460 254.800 ;
      RECT 77.420 1.400 77.700 254.800 ;
      RECT 79.660 1.400 79.940 254.800 ;
      RECT 81.900 1.400 82.180 254.800 ;
      RECT 84.140 1.400 84.420 254.800 ;
      RECT 86.380 1.400 86.660 254.800 ;
      RECT 88.620 1.400 88.900 254.800 ;
      RECT 90.860 1.400 91.140 254.800 ;
      RECT 93.100 1.400 93.380 254.800 ;
      RECT 95.340 1.400 95.620 254.800 ;
      RECT 97.580 1.400 97.860 254.800 ;
      RECT 99.820 1.400 100.100 254.800 ;
      RECT 102.060 1.400 102.340 254.800 ;
      RECT 104.300 1.400 104.580 254.800 ;
      RECT 106.540 1.400 106.820 254.800 ;
      RECT 108.780 1.400 109.060 254.800 ;
      RECT 111.020 1.400 111.300 254.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 254.800 ;
      RECT 4.620 1.400 4.900 254.800 ;
      RECT 6.860 1.400 7.140 254.800 ;
      RECT 9.100 1.400 9.380 254.800 ;
      RECT 11.340 1.400 11.620 254.800 ;
      RECT 13.580 1.400 13.860 254.800 ;
      RECT 15.820 1.400 16.100 254.800 ;
      RECT 18.060 1.400 18.340 254.800 ;
      RECT 20.300 1.400 20.580 254.800 ;
      RECT 22.540 1.400 22.820 254.800 ;
      RECT 24.780 1.400 25.060 254.800 ;
      RECT 27.020 1.400 27.300 254.800 ;
      RECT 29.260 1.400 29.540 254.800 ;
      RECT 31.500 1.400 31.780 254.800 ;
      RECT 33.740 1.400 34.020 254.800 ;
      RECT 35.980 1.400 36.260 254.800 ;
      RECT 38.220 1.400 38.500 254.800 ;
      RECT 40.460 1.400 40.740 254.800 ;
      RECT 42.700 1.400 42.980 254.800 ;
      RECT 44.940 1.400 45.220 254.800 ;
      RECT 47.180 1.400 47.460 254.800 ;
      RECT 49.420 1.400 49.700 254.800 ;
      RECT 51.660 1.400 51.940 254.800 ;
      RECT 53.900 1.400 54.180 254.800 ;
      RECT 56.140 1.400 56.420 254.800 ;
      RECT 58.380 1.400 58.660 254.800 ;
      RECT 60.620 1.400 60.900 254.800 ;
      RECT 62.860 1.400 63.140 254.800 ;
      RECT 65.100 1.400 65.380 254.800 ;
      RECT 67.340 1.400 67.620 254.800 ;
      RECT 69.580 1.400 69.860 254.800 ;
      RECT 71.820 1.400 72.100 254.800 ;
      RECT 74.060 1.400 74.340 254.800 ;
      RECT 76.300 1.400 76.580 254.800 ;
      RECT 78.540 1.400 78.820 254.800 ;
      RECT 80.780 1.400 81.060 254.800 ;
      RECT 83.020 1.400 83.300 254.800 ;
      RECT 85.260 1.400 85.540 254.800 ;
      RECT 87.500 1.400 87.780 254.800 ;
      RECT 89.740 1.400 90.020 254.800 ;
      RECT 91.980 1.400 92.260 254.800 ;
      RECT 94.220 1.400 94.500 254.800 ;
      RECT 96.460 1.400 96.740 254.800 ;
      RECT 98.700 1.400 98.980 254.800 ;
      RECT 100.940 1.400 101.220 254.800 ;
      RECT 103.180 1.400 103.460 254.800 ;
      RECT 105.420 1.400 105.700 254.800 ;
      RECT 107.660 1.400 107.940 254.800 ;
      RECT 109.900 1.400 110.180 254.800 ;
      RECT 112.140 1.400 112.420 254.800 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 114.000 256.200 ;
    LAYER metal2 ;
    RECT 0 0 114.000 256.200 ;
    LAYER metal3 ;
    RECT 0.070 0 114.000 256.200 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 3.465 ;
    RECT 0 3.535 0.070 5.565 ;
    RECT 0 5.635 0.070 7.665 ;
    RECT 0 7.735 0.070 9.765 ;
    RECT 0 9.835 0.070 11.865 ;
    RECT 0 11.935 0.070 13.965 ;
    RECT 0 14.035 0.070 16.065 ;
    RECT 0 16.135 0.070 18.165 ;
    RECT 0 18.235 0.070 20.265 ;
    RECT 0 20.335 0.070 22.365 ;
    RECT 0 22.435 0.070 24.465 ;
    RECT 0 24.535 0.070 26.565 ;
    RECT 0 26.635 0.070 28.665 ;
    RECT 0 28.735 0.070 30.765 ;
    RECT 0 30.835 0.070 32.865 ;
    RECT 0 32.935 0.070 34.965 ;
    RECT 0 35.035 0.070 37.065 ;
    RECT 0 37.135 0.070 39.165 ;
    RECT 0 39.235 0.070 41.265 ;
    RECT 0 41.335 0.070 43.365 ;
    RECT 0 43.435 0.070 45.465 ;
    RECT 0 45.535 0.070 47.565 ;
    RECT 0 47.635 0.070 49.665 ;
    RECT 0 49.735 0.070 51.765 ;
    RECT 0 51.835 0.070 53.865 ;
    RECT 0 53.935 0.070 55.965 ;
    RECT 0 56.035 0.070 58.065 ;
    RECT 0 58.135 0.070 60.165 ;
    RECT 0 60.235 0.070 62.265 ;
    RECT 0 62.335 0.070 64.365 ;
    RECT 0 64.435 0.070 66.465 ;
    RECT 0 66.535 0.070 66.605 ;
    RECT 0 66.675 0.070 68.705 ;
    RECT 0 68.775 0.070 70.805 ;
    RECT 0 70.875 0.070 72.905 ;
    RECT 0 72.975 0.070 75.005 ;
    RECT 0 75.075 0.070 77.105 ;
    RECT 0 77.175 0.070 79.205 ;
    RECT 0 79.275 0.070 81.305 ;
    RECT 0 81.375 0.070 83.405 ;
    RECT 0 83.475 0.070 85.505 ;
    RECT 0 85.575 0.070 87.605 ;
    RECT 0 87.675 0.070 89.705 ;
    RECT 0 89.775 0.070 91.805 ;
    RECT 0 91.875 0.070 93.905 ;
    RECT 0 93.975 0.070 96.005 ;
    RECT 0 96.075 0.070 98.105 ;
    RECT 0 98.175 0.070 100.205 ;
    RECT 0 100.275 0.070 102.305 ;
    RECT 0 102.375 0.070 104.405 ;
    RECT 0 104.475 0.070 106.505 ;
    RECT 0 106.575 0.070 108.605 ;
    RECT 0 108.675 0.070 110.705 ;
    RECT 0 110.775 0.070 112.805 ;
    RECT 0 112.875 0.070 114.905 ;
    RECT 0 114.975 0.070 117.005 ;
    RECT 0 117.075 0.070 119.105 ;
    RECT 0 119.175 0.070 121.205 ;
    RECT 0 121.275 0.070 123.305 ;
    RECT 0 123.375 0.070 125.405 ;
    RECT 0 125.475 0.070 127.505 ;
    RECT 0 127.575 0.070 129.605 ;
    RECT 0 129.675 0.070 131.705 ;
    RECT 0 131.775 0.070 131.845 ;
    RECT 0 131.915 0.070 133.945 ;
    RECT 0 134.015 0.070 136.045 ;
    RECT 0 136.115 0.070 138.145 ;
    RECT 0 138.215 0.070 140.245 ;
    RECT 0 140.315 0.070 142.345 ;
    RECT 0 142.415 0.070 144.445 ;
    RECT 0 144.515 0.070 146.545 ;
    RECT 0 146.615 0.070 148.645 ;
    RECT 0 148.715 0.070 150.745 ;
    RECT 0 150.815 0.070 152.845 ;
    RECT 0 152.915 0.070 154.945 ;
    RECT 0 155.015 0.070 157.045 ;
    RECT 0 157.115 0.070 159.145 ;
    RECT 0 159.215 0.070 161.245 ;
    RECT 0 161.315 0.070 163.345 ;
    RECT 0 163.415 0.070 165.445 ;
    RECT 0 165.515 0.070 167.545 ;
    RECT 0 167.615 0.070 169.645 ;
    RECT 0 169.715 0.070 171.745 ;
    RECT 0 171.815 0.070 173.845 ;
    RECT 0 173.915 0.070 175.945 ;
    RECT 0 176.015 0.070 178.045 ;
    RECT 0 178.115 0.070 180.145 ;
    RECT 0 180.215 0.070 182.245 ;
    RECT 0 182.315 0.070 184.345 ;
    RECT 0 184.415 0.070 186.445 ;
    RECT 0 186.515 0.070 188.545 ;
    RECT 0 188.615 0.070 190.645 ;
    RECT 0 190.715 0.070 192.745 ;
    RECT 0 192.815 0.070 194.845 ;
    RECT 0 194.915 0.070 196.945 ;
    RECT 0 197.015 0.070 197.085 ;
    RECT 0 197.155 0.070 199.185 ;
    RECT 0 199.255 0.070 201.285 ;
    RECT 0 201.355 0.070 203.385 ;
    RECT 0 203.455 0.070 205.485 ;
    RECT 0 205.555 0.070 207.585 ;
    RECT 0 207.655 0.070 209.685 ;
    RECT 0 209.755 0.070 211.785 ;
    RECT 0 211.855 0.070 213.885 ;
    RECT 0 213.955 0.070 214.025 ;
    RECT 0 214.095 0.070 216.125 ;
    RECT 0 216.195 0.070 218.225 ;
    RECT 0 218.295 0.070 256.200 ;
    LAYER metal4 ;
    RECT 0 0 114.000 1.400 ;
    RECT 0 254.800 114.000 256.200 ;
    RECT 0.000 1.400 1.260 254.800 ;
    RECT 1.540 1.400 2.380 254.800 ;
    RECT 2.660 1.400 3.500 254.800 ;
    RECT 3.780 1.400 4.620 254.800 ;
    RECT 4.900 1.400 5.740 254.800 ;
    RECT 6.020 1.400 6.860 254.800 ;
    RECT 7.140 1.400 7.980 254.800 ;
    RECT 8.260 1.400 9.100 254.800 ;
    RECT 9.380 1.400 10.220 254.800 ;
    RECT 10.500 1.400 11.340 254.800 ;
    RECT 11.620 1.400 12.460 254.800 ;
    RECT 12.740 1.400 13.580 254.800 ;
    RECT 13.860 1.400 14.700 254.800 ;
    RECT 14.980 1.400 15.820 254.800 ;
    RECT 16.100 1.400 16.940 254.800 ;
    RECT 17.220 1.400 18.060 254.800 ;
    RECT 18.340 1.400 19.180 254.800 ;
    RECT 19.460 1.400 20.300 254.800 ;
    RECT 20.580 1.400 21.420 254.800 ;
    RECT 21.700 1.400 22.540 254.800 ;
    RECT 22.820 1.400 23.660 254.800 ;
    RECT 23.940 1.400 24.780 254.800 ;
    RECT 25.060 1.400 25.900 254.800 ;
    RECT 26.180 1.400 27.020 254.800 ;
    RECT 27.300 1.400 28.140 254.800 ;
    RECT 28.420 1.400 29.260 254.800 ;
    RECT 29.540 1.400 30.380 254.800 ;
    RECT 30.660 1.400 31.500 254.800 ;
    RECT 31.780 1.400 32.620 254.800 ;
    RECT 32.900 1.400 33.740 254.800 ;
    RECT 34.020 1.400 34.860 254.800 ;
    RECT 35.140 1.400 35.980 254.800 ;
    RECT 36.260 1.400 37.100 254.800 ;
    RECT 37.380 1.400 38.220 254.800 ;
    RECT 38.500 1.400 39.340 254.800 ;
    RECT 39.620 1.400 40.460 254.800 ;
    RECT 40.740 1.400 41.580 254.800 ;
    RECT 41.860 1.400 42.700 254.800 ;
    RECT 42.980 1.400 43.820 254.800 ;
    RECT 44.100 1.400 44.940 254.800 ;
    RECT 45.220 1.400 46.060 254.800 ;
    RECT 46.340 1.400 47.180 254.800 ;
    RECT 47.460 1.400 48.300 254.800 ;
    RECT 48.580 1.400 49.420 254.800 ;
    RECT 49.700 1.400 50.540 254.800 ;
    RECT 50.820 1.400 51.660 254.800 ;
    RECT 51.940 1.400 52.780 254.800 ;
    RECT 53.060 1.400 53.900 254.800 ;
    RECT 54.180 1.400 55.020 254.800 ;
    RECT 55.300 1.400 56.140 254.800 ;
    RECT 56.420 1.400 57.260 254.800 ;
    RECT 57.540 1.400 58.380 254.800 ;
    RECT 58.660 1.400 59.500 254.800 ;
    RECT 59.780 1.400 60.620 254.800 ;
    RECT 60.900 1.400 61.740 254.800 ;
    RECT 62.020 1.400 62.860 254.800 ;
    RECT 63.140 1.400 63.980 254.800 ;
    RECT 64.260 1.400 65.100 254.800 ;
    RECT 65.380 1.400 66.220 254.800 ;
    RECT 66.500 1.400 67.340 254.800 ;
    RECT 67.620 1.400 68.460 254.800 ;
    RECT 68.740 1.400 69.580 254.800 ;
    RECT 69.860 1.400 70.700 254.800 ;
    RECT 70.980 1.400 71.820 254.800 ;
    RECT 72.100 1.400 72.940 254.800 ;
    RECT 73.220 1.400 74.060 254.800 ;
    RECT 74.340 1.400 75.180 254.800 ;
    RECT 75.460 1.400 76.300 254.800 ;
    RECT 76.580 1.400 77.420 254.800 ;
    RECT 77.700 1.400 78.540 254.800 ;
    RECT 78.820 1.400 79.660 254.800 ;
    RECT 79.940 1.400 80.780 254.800 ;
    RECT 81.060 1.400 81.900 254.800 ;
    RECT 82.180 1.400 83.020 254.800 ;
    RECT 83.300 1.400 84.140 254.800 ;
    RECT 84.420 1.400 85.260 254.800 ;
    RECT 85.540 1.400 86.380 254.800 ;
    RECT 86.660 1.400 87.500 254.800 ;
    RECT 87.780 1.400 88.620 254.800 ;
    RECT 88.900 1.400 89.740 254.800 ;
    RECT 90.020 1.400 90.860 254.800 ;
    RECT 91.140 1.400 91.980 254.800 ;
    RECT 92.260 1.400 93.100 254.800 ;
    RECT 93.380 1.400 94.220 254.800 ;
    RECT 94.500 1.400 95.340 254.800 ;
    RECT 95.620 1.400 96.460 254.800 ;
    RECT 96.740 1.400 97.580 254.800 ;
    RECT 97.860 1.400 98.700 254.800 ;
    RECT 98.980 1.400 99.820 254.800 ;
    RECT 100.100 1.400 100.940 254.800 ;
    RECT 101.220 1.400 102.060 254.800 ;
    RECT 102.340 1.400 103.180 254.800 ;
    RECT 103.460 1.400 104.300 254.800 ;
    RECT 104.580 1.400 105.420 254.800 ;
    RECT 105.700 1.400 106.540 254.800 ;
    RECT 106.820 1.400 107.660 254.800 ;
    RECT 107.940 1.400 108.780 254.800 ;
    RECT 109.060 1.400 109.900 254.800 ;
    RECT 110.180 1.400 111.020 254.800 ;
    RECT 111.300 1.400 112.140 254.800 ;
    RECT 112.420 1.400 114.000 254.800 ;
    LAYER OVERLAP ;
    RECT 0 0 114.000 256.200 ;
  END
END liteeth_1rw1r_32w384d_8_sram

END LIBRARY
