VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_512x256_1r1w
  FOREIGN fakeram_512x256_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 1302.720 BY 1569.440 ;
  CLASS BLOCK ;
  PIN w0_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 6.650 0.800 6.950 ;
    END
  END w0_mask_in[0]
  PIN w0_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 8.010 0.800 8.310 ;
    END
  END w0_mask_in[1]
  PIN w0_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 9.370 0.800 9.670 ;
    END
  END w0_mask_in[2]
  PIN w0_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 10.730 0.800 11.030 ;
    END
  END w0_mask_in[3]
  PIN w0_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 12.090 0.800 12.390 ;
    END
  END w0_mask_in[4]
  PIN w0_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 13.450 0.800 13.750 ;
    END
  END w0_mask_in[5]
  PIN w0_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.810 0.800 15.110 ;
    END
  END w0_mask_in[6]
  PIN w0_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 16.170 0.800 16.470 ;
    END
  END w0_mask_in[7]
  PIN w0_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 17.530 0.800 17.830 ;
    END
  END w0_mask_in[8]
  PIN w0_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 18.890 0.800 19.190 ;
    END
  END w0_mask_in[9]
  PIN w0_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.250 0.800 20.550 ;
    END
  END w0_mask_in[10]
  PIN w0_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 21.610 0.800 21.910 ;
    END
  END w0_mask_in[11]
  PIN w0_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.970 0.800 23.270 ;
    END
  END w0_mask_in[12]
  PIN w0_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 24.330 0.800 24.630 ;
    END
  END w0_mask_in[13]
  PIN w0_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 25.690 0.800 25.990 ;
    END
  END w0_mask_in[14]
  PIN w0_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 27.050 0.800 27.350 ;
    END
  END w0_mask_in[15]
  PIN w0_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 28.410 0.800 28.710 ;
    END
  END w0_mask_in[16]
  PIN w0_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 29.770 0.800 30.070 ;
    END
  END w0_mask_in[17]
  PIN w0_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.130 0.800 31.430 ;
    END
  END w0_mask_in[18]
  PIN w0_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 32.490 0.800 32.790 ;
    END
  END w0_mask_in[19]
  PIN w0_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 33.850 0.800 34.150 ;
    END
  END w0_mask_in[20]
  PIN w0_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 35.210 0.800 35.510 ;
    END
  END w0_mask_in[21]
  PIN w0_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 36.570 0.800 36.870 ;
    END
  END w0_mask_in[22]
  PIN w0_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.930 0.800 38.230 ;
    END
  END w0_mask_in[23]
  PIN w0_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.290 0.800 39.590 ;
    END
  END w0_mask_in[24]
  PIN w0_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.650 0.800 40.950 ;
    END
  END w0_mask_in[25]
  PIN w0_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 42.010 0.800 42.310 ;
    END
  END w0_mask_in[26]
  PIN w0_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 43.370 0.800 43.670 ;
    END
  END w0_mask_in[27]
  PIN w0_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 44.730 0.800 45.030 ;
    END
  END w0_mask_in[28]
  PIN w0_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 46.090 0.800 46.390 ;
    END
  END w0_mask_in[29]
  PIN w0_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 47.450 0.800 47.750 ;
    END
  END w0_mask_in[30]
  PIN w0_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 48.810 0.800 49.110 ;
    END
  END w0_mask_in[31]
  PIN w0_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 50.170 0.800 50.470 ;
    END
  END w0_mask_in[32]
  PIN w0_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 51.530 0.800 51.830 ;
    END
  END w0_mask_in[33]
  PIN w0_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 52.890 0.800 53.190 ;
    END
  END w0_mask_in[34]
  PIN w0_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 54.250 0.800 54.550 ;
    END
  END w0_mask_in[35]
  PIN w0_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.610 0.800 55.910 ;
    END
  END w0_mask_in[36]
  PIN w0_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 56.970 0.800 57.270 ;
    END
  END w0_mask_in[37]
  PIN w0_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 58.330 0.800 58.630 ;
    END
  END w0_mask_in[38]
  PIN w0_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 59.690 0.800 59.990 ;
    END
  END w0_mask_in[39]
  PIN w0_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 61.050 0.800 61.350 ;
    END
  END w0_mask_in[40]
  PIN w0_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 62.410 0.800 62.710 ;
    END
  END w0_mask_in[41]
  PIN w0_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 63.770 0.800 64.070 ;
    END
  END w0_mask_in[42]
  PIN w0_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 65.130 0.800 65.430 ;
    END
  END w0_mask_in[43]
  PIN w0_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 66.490 0.800 66.790 ;
    END
  END w0_mask_in[44]
  PIN w0_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.850 0.800 68.150 ;
    END
  END w0_mask_in[45]
  PIN w0_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 69.210 0.800 69.510 ;
    END
  END w0_mask_in[46]
  PIN w0_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 70.570 0.800 70.870 ;
    END
  END w0_mask_in[47]
  PIN w0_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.930 0.800 72.230 ;
    END
  END w0_mask_in[48]
  PIN w0_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 73.290 0.800 73.590 ;
    END
  END w0_mask_in[49]
  PIN w0_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 74.650 0.800 74.950 ;
    END
  END w0_mask_in[50]
  PIN w0_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.010 0.800 76.310 ;
    END
  END w0_mask_in[51]
  PIN w0_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 77.370 0.800 77.670 ;
    END
  END w0_mask_in[52]
  PIN w0_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 78.730 0.800 79.030 ;
    END
  END w0_mask_in[53]
  PIN w0_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 80.090 0.800 80.390 ;
    END
  END w0_mask_in[54]
  PIN w0_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 81.450 0.800 81.750 ;
    END
  END w0_mask_in[55]
  PIN w0_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 82.810 0.800 83.110 ;
    END
  END w0_mask_in[56]
  PIN w0_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 84.170 0.800 84.470 ;
    END
  END w0_mask_in[57]
  PIN w0_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 85.530 0.800 85.830 ;
    END
  END w0_mask_in[58]
  PIN w0_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 86.890 0.800 87.190 ;
    END
  END w0_mask_in[59]
  PIN w0_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 88.250 0.800 88.550 ;
    END
  END w0_mask_in[60]
  PIN w0_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.610 0.800 89.910 ;
    END
  END w0_mask_in[61]
  PIN w0_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 90.970 0.800 91.270 ;
    END
  END w0_mask_in[62]
  PIN w0_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 92.330 0.800 92.630 ;
    END
  END w0_mask_in[63]
  PIN w0_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 93.690 0.800 93.990 ;
    END
  END w0_mask_in[64]
  PIN w0_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 95.050 0.800 95.350 ;
    END
  END w0_mask_in[65]
  PIN w0_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 96.410 0.800 96.710 ;
    END
  END w0_mask_in[66]
  PIN w0_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 97.770 0.800 98.070 ;
    END
  END w0_mask_in[67]
  PIN w0_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 99.130 0.800 99.430 ;
    END
  END w0_mask_in[68]
  PIN w0_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 100.490 0.800 100.790 ;
    END
  END w0_mask_in[69]
  PIN w0_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 101.850 0.800 102.150 ;
    END
  END w0_mask_in[70]
  PIN w0_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 103.210 0.800 103.510 ;
    END
  END w0_mask_in[71]
  PIN w0_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 104.570 0.800 104.870 ;
    END
  END w0_mask_in[72]
  PIN w0_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 105.930 0.800 106.230 ;
    END
  END w0_mask_in[73]
  PIN w0_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 107.290 0.800 107.590 ;
    END
  END w0_mask_in[74]
  PIN w0_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 108.650 0.800 108.950 ;
    END
  END w0_mask_in[75]
  PIN w0_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 110.010 0.800 110.310 ;
    END
  END w0_mask_in[76]
  PIN w0_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 111.370 0.800 111.670 ;
    END
  END w0_mask_in[77]
  PIN w0_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 112.730 0.800 113.030 ;
    END
  END w0_mask_in[78]
  PIN w0_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 114.090 0.800 114.390 ;
    END
  END w0_mask_in[79]
  PIN w0_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 115.450 0.800 115.750 ;
    END
  END w0_mask_in[80]
  PIN w0_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 116.810 0.800 117.110 ;
    END
  END w0_mask_in[81]
  PIN w0_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 118.170 0.800 118.470 ;
    END
  END w0_mask_in[82]
  PIN w0_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 119.530 0.800 119.830 ;
    END
  END w0_mask_in[83]
  PIN w0_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 120.890 0.800 121.190 ;
    END
  END w0_mask_in[84]
  PIN w0_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 122.250 0.800 122.550 ;
    END
  END w0_mask_in[85]
  PIN w0_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 123.610 0.800 123.910 ;
    END
  END w0_mask_in[86]
  PIN w0_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 124.970 0.800 125.270 ;
    END
  END w0_mask_in[87]
  PIN w0_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 126.330 0.800 126.630 ;
    END
  END w0_mask_in[88]
  PIN w0_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 127.690 0.800 127.990 ;
    END
  END w0_mask_in[89]
  PIN w0_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 129.050 0.800 129.350 ;
    END
  END w0_mask_in[90]
  PIN w0_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 130.410 0.800 130.710 ;
    END
  END w0_mask_in[91]
  PIN w0_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 131.770 0.800 132.070 ;
    END
  END w0_mask_in[92]
  PIN w0_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 133.130 0.800 133.430 ;
    END
  END w0_mask_in[93]
  PIN w0_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 134.490 0.800 134.790 ;
    END
  END w0_mask_in[94]
  PIN w0_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 135.850 0.800 136.150 ;
    END
  END w0_mask_in[95]
  PIN w0_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 137.210 0.800 137.510 ;
    END
  END w0_mask_in[96]
  PIN w0_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 138.570 0.800 138.870 ;
    END
  END w0_mask_in[97]
  PIN w0_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.930 0.800 140.230 ;
    END
  END w0_mask_in[98]
  PIN w0_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 141.290 0.800 141.590 ;
    END
  END w0_mask_in[99]
  PIN w0_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 142.650 0.800 142.950 ;
    END
  END w0_mask_in[100]
  PIN w0_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 144.010 0.800 144.310 ;
    END
  END w0_mask_in[101]
  PIN w0_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 145.370 0.800 145.670 ;
    END
  END w0_mask_in[102]
  PIN w0_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 146.730 0.800 147.030 ;
    END
  END w0_mask_in[103]
  PIN w0_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 148.090 0.800 148.390 ;
    END
  END w0_mask_in[104]
  PIN w0_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 149.450 0.800 149.750 ;
    END
  END w0_mask_in[105]
  PIN w0_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 150.810 0.800 151.110 ;
    END
  END w0_mask_in[106]
  PIN w0_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 152.170 0.800 152.470 ;
    END
  END w0_mask_in[107]
  PIN w0_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 153.530 0.800 153.830 ;
    END
  END w0_mask_in[108]
  PIN w0_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 154.890 0.800 155.190 ;
    END
  END w0_mask_in[109]
  PIN w0_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 156.250 0.800 156.550 ;
    END
  END w0_mask_in[110]
  PIN w0_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 157.610 0.800 157.910 ;
    END
  END w0_mask_in[111]
  PIN w0_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 158.970 0.800 159.270 ;
    END
  END w0_mask_in[112]
  PIN w0_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 160.330 0.800 160.630 ;
    END
  END w0_mask_in[113]
  PIN w0_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 161.690 0.800 161.990 ;
    END
  END w0_mask_in[114]
  PIN w0_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 163.050 0.800 163.350 ;
    END
  END w0_mask_in[115]
  PIN w0_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 164.410 0.800 164.710 ;
    END
  END w0_mask_in[116]
  PIN w0_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 165.770 0.800 166.070 ;
    END
  END w0_mask_in[117]
  PIN w0_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 167.130 0.800 167.430 ;
    END
  END w0_mask_in[118]
  PIN w0_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 168.490 0.800 168.790 ;
    END
  END w0_mask_in[119]
  PIN w0_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 169.850 0.800 170.150 ;
    END
  END w0_mask_in[120]
  PIN w0_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 171.210 0.800 171.510 ;
    END
  END w0_mask_in[121]
  PIN w0_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 172.570 0.800 172.870 ;
    END
  END w0_mask_in[122]
  PIN w0_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 173.930 0.800 174.230 ;
    END
  END w0_mask_in[123]
  PIN w0_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 175.290 0.800 175.590 ;
    END
  END w0_mask_in[124]
  PIN w0_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 176.650 0.800 176.950 ;
    END
  END w0_mask_in[125]
  PIN w0_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 178.010 0.800 178.310 ;
    END
  END w0_mask_in[126]
  PIN w0_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 179.370 0.800 179.670 ;
    END
  END w0_mask_in[127]
  PIN w0_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 180.730 0.800 181.030 ;
    END
  END w0_mask_in[128]
  PIN w0_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 182.090 0.800 182.390 ;
    END
  END w0_mask_in[129]
  PIN w0_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 183.450 0.800 183.750 ;
    END
  END w0_mask_in[130]
  PIN w0_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 184.810 0.800 185.110 ;
    END
  END w0_mask_in[131]
  PIN w0_mask_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 186.170 0.800 186.470 ;
    END
  END w0_mask_in[132]
  PIN w0_mask_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 187.530 0.800 187.830 ;
    END
  END w0_mask_in[133]
  PIN w0_mask_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 188.890 0.800 189.190 ;
    END
  END w0_mask_in[134]
  PIN w0_mask_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 190.250 0.800 190.550 ;
    END
  END w0_mask_in[135]
  PIN w0_mask_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 191.610 0.800 191.910 ;
    END
  END w0_mask_in[136]
  PIN w0_mask_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 192.970 0.800 193.270 ;
    END
  END w0_mask_in[137]
  PIN w0_mask_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 194.330 0.800 194.630 ;
    END
  END w0_mask_in[138]
  PIN w0_mask_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 195.690 0.800 195.990 ;
    END
  END w0_mask_in[139]
  PIN w0_mask_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 197.050 0.800 197.350 ;
    END
  END w0_mask_in[140]
  PIN w0_mask_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 198.410 0.800 198.710 ;
    END
  END w0_mask_in[141]
  PIN w0_mask_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 199.770 0.800 200.070 ;
    END
  END w0_mask_in[142]
  PIN w0_mask_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 201.130 0.800 201.430 ;
    END
  END w0_mask_in[143]
  PIN w0_mask_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 202.490 0.800 202.790 ;
    END
  END w0_mask_in[144]
  PIN w0_mask_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 203.850 0.800 204.150 ;
    END
  END w0_mask_in[145]
  PIN w0_mask_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 205.210 0.800 205.510 ;
    END
  END w0_mask_in[146]
  PIN w0_mask_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 206.570 0.800 206.870 ;
    END
  END w0_mask_in[147]
  PIN w0_mask_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 207.930 0.800 208.230 ;
    END
  END w0_mask_in[148]
  PIN w0_mask_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 209.290 0.800 209.590 ;
    END
  END w0_mask_in[149]
  PIN w0_mask_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 210.650 0.800 210.950 ;
    END
  END w0_mask_in[150]
  PIN w0_mask_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 212.010 0.800 212.310 ;
    END
  END w0_mask_in[151]
  PIN w0_mask_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 213.370 0.800 213.670 ;
    END
  END w0_mask_in[152]
  PIN w0_mask_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 214.730 0.800 215.030 ;
    END
  END w0_mask_in[153]
  PIN w0_mask_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 216.090 0.800 216.390 ;
    END
  END w0_mask_in[154]
  PIN w0_mask_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 217.450 0.800 217.750 ;
    END
  END w0_mask_in[155]
  PIN w0_mask_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 218.810 0.800 219.110 ;
    END
  END w0_mask_in[156]
  PIN w0_mask_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 220.170 0.800 220.470 ;
    END
  END w0_mask_in[157]
  PIN w0_mask_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 221.530 0.800 221.830 ;
    END
  END w0_mask_in[158]
  PIN w0_mask_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 222.890 0.800 223.190 ;
    END
  END w0_mask_in[159]
  PIN w0_mask_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 224.250 0.800 224.550 ;
    END
  END w0_mask_in[160]
  PIN w0_mask_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 225.610 0.800 225.910 ;
    END
  END w0_mask_in[161]
  PIN w0_mask_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 226.970 0.800 227.270 ;
    END
  END w0_mask_in[162]
  PIN w0_mask_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 228.330 0.800 228.630 ;
    END
  END w0_mask_in[163]
  PIN w0_mask_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 229.690 0.800 229.990 ;
    END
  END w0_mask_in[164]
  PIN w0_mask_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 231.050 0.800 231.350 ;
    END
  END w0_mask_in[165]
  PIN w0_mask_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 232.410 0.800 232.710 ;
    END
  END w0_mask_in[166]
  PIN w0_mask_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 233.770 0.800 234.070 ;
    END
  END w0_mask_in[167]
  PIN w0_mask_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 235.130 0.800 235.430 ;
    END
  END w0_mask_in[168]
  PIN w0_mask_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 236.490 0.800 236.790 ;
    END
  END w0_mask_in[169]
  PIN w0_mask_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 237.850 0.800 238.150 ;
    END
  END w0_mask_in[170]
  PIN w0_mask_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 239.210 0.800 239.510 ;
    END
  END w0_mask_in[171]
  PIN w0_mask_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 240.570 0.800 240.870 ;
    END
  END w0_mask_in[172]
  PIN w0_mask_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 241.930 0.800 242.230 ;
    END
  END w0_mask_in[173]
  PIN w0_mask_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 243.290 0.800 243.590 ;
    END
  END w0_mask_in[174]
  PIN w0_mask_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 244.650 0.800 244.950 ;
    END
  END w0_mask_in[175]
  PIN w0_mask_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 246.010 0.800 246.310 ;
    END
  END w0_mask_in[176]
  PIN w0_mask_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 247.370 0.800 247.670 ;
    END
  END w0_mask_in[177]
  PIN w0_mask_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 248.730 0.800 249.030 ;
    END
  END w0_mask_in[178]
  PIN w0_mask_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 250.090 0.800 250.390 ;
    END
  END w0_mask_in[179]
  PIN w0_mask_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 251.450 0.800 251.750 ;
    END
  END w0_mask_in[180]
  PIN w0_mask_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 252.810 0.800 253.110 ;
    END
  END w0_mask_in[181]
  PIN w0_mask_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 254.170 0.800 254.470 ;
    END
  END w0_mask_in[182]
  PIN w0_mask_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 255.530 0.800 255.830 ;
    END
  END w0_mask_in[183]
  PIN w0_mask_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 256.890 0.800 257.190 ;
    END
  END w0_mask_in[184]
  PIN w0_mask_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 258.250 0.800 258.550 ;
    END
  END w0_mask_in[185]
  PIN w0_mask_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 259.610 0.800 259.910 ;
    END
  END w0_mask_in[186]
  PIN w0_mask_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 260.970 0.800 261.270 ;
    END
  END w0_mask_in[187]
  PIN w0_mask_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 262.330 0.800 262.630 ;
    END
  END w0_mask_in[188]
  PIN w0_mask_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 263.690 0.800 263.990 ;
    END
  END w0_mask_in[189]
  PIN w0_mask_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 265.050 0.800 265.350 ;
    END
  END w0_mask_in[190]
  PIN w0_mask_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 266.410 0.800 266.710 ;
    END
  END w0_mask_in[191]
  PIN w0_mask_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 267.770 0.800 268.070 ;
    END
  END w0_mask_in[192]
  PIN w0_mask_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 269.130 0.800 269.430 ;
    END
  END w0_mask_in[193]
  PIN w0_mask_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 270.490 0.800 270.790 ;
    END
  END w0_mask_in[194]
  PIN w0_mask_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 271.850 0.800 272.150 ;
    END
  END w0_mask_in[195]
  PIN w0_mask_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 273.210 0.800 273.510 ;
    END
  END w0_mask_in[196]
  PIN w0_mask_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 274.570 0.800 274.870 ;
    END
  END w0_mask_in[197]
  PIN w0_mask_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 275.930 0.800 276.230 ;
    END
  END w0_mask_in[198]
  PIN w0_mask_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 277.290 0.800 277.590 ;
    END
  END w0_mask_in[199]
  PIN w0_mask_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 278.650 0.800 278.950 ;
    END
  END w0_mask_in[200]
  PIN w0_mask_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 280.010 0.800 280.310 ;
    END
  END w0_mask_in[201]
  PIN w0_mask_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 281.370 0.800 281.670 ;
    END
  END w0_mask_in[202]
  PIN w0_mask_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 282.730 0.800 283.030 ;
    END
  END w0_mask_in[203]
  PIN w0_mask_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 284.090 0.800 284.390 ;
    END
  END w0_mask_in[204]
  PIN w0_mask_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 285.450 0.800 285.750 ;
    END
  END w0_mask_in[205]
  PIN w0_mask_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 286.810 0.800 287.110 ;
    END
  END w0_mask_in[206]
  PIN w0_mask_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 288.170 0.800 288.470 ;
    END
  END w0_mask_in[207]
  PIN w0_mask_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 289.530 0.800 289.830 ;
    END
  END w0_mask_in[208]
  PIN w0_mask_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 290.890 0.800 291.190 ;
    END
  END w0_mask_in[209]
  PIN w0_mask_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 292.250 0.800 292.550 ;
    END
  END w0_mask_in[210]
  PIN w0_mask_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 293.610 0.800 293.910 ;
    END
  END w0_mask_in[211]
  PIN w0_mask_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 294.970 0.800 295.270 ;
    END
  END w0_mask_in[212]
  PIN w0_mask_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 296.330 0.800 296.630 ;
    END
  END w0_mask_in[213]
  PIN w0_mask_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 297.690 0.800 297.990 ;
    END
  END w0_mask_in[214]
  PIN w0_mask_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 299.050 0.800 299.350 ;
    END
  END w0_mask_in[215]
  PIN w0_mask_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 300.410 0.800 300.710 ;
    END
  END w0_mask_in[216]
  PIN w0_mask_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 301.770 0.800 302.070 ;
    END
  END w0_mask_in[217]
  PIN w0_mask_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 303.130 0.800 303.430 ;
    END
  END w0_mask_in[218]
  PIN w0_mask_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 304.490 0.800 304.790 ;
    END
  END w0_mask_in[219]
  PIN w0_mask_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 305.850 0.800 306.150 ;
    END
  END w0_mask_in[220]
  PIN w0_mask_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 307.210 0.800 307.510 ;
    END
  END w0_mask_in[221]
  PIN w0_mask_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 308.570 0.800 308.870 ;
    END
  END w0_mask_in[222]
  PIN w0_mask_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 309.930 0.800 310.230 ;
    END
  END w0_mask_in[223]
  PIN w0_mask_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 311.290 0.800 311.590 ;
    END
  END w0_mask_in[224]
  PIN w0_mask_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 312.650 0.800 312.950 ;
    END
  END w0_mask_in[225]
  PIN w0_mask_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 314.010 0.800 314.310 ;
    END
  END w0_mask_in[226]
  PIN w0_mask_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 315.370 0.800 315.670 ;
    END
  END w0_mask_in[227]
  PIN w0_mask_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 316.730 0.800 317.030 ;
    END
  END w0_mask_in[228]
  PIN w0_mask_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 318.090 0.800 318.390 ;
    END
  END w0_mask_in[229]
  PIN w0_mask_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 319.450 0.800 319.750 ;
    END
  END w0_mask_in[230]
  PIN w0_mask_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 320.810 0.800 321.110 ;
    END
  END w0_mask_in[231]
  PIN w0_mask_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 322.170 0.800 322.470 ;
    END
  END w0_mask_in[232]
  PIN w0_mask_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 323.530 0.800 323.830 ;
    END
  END w0_mask_in[233]
  PIN w0_mask_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 324.890 0.800 325.190 ;
    END
  END w0_mask_in[234]
  PIN w0_mask_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 326.250 0.800 326.550 ;
    END
  END w0_mask_in[235]
  PIN w0_mask_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 327.610 0.800 327.910 ;
    END
  END w0_mask_in[236]
  PIN w0_mask_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 328.970 0.800 329.270 ;
    END
  END w0_mask_in[237]
  PIN w0_mask_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 330.330 0.800 330.630 ;
    END
  END w0_mask_in[238]
  PIN w0_mask_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 331.690 0.800 331.990 ;
    END
  END w0_mask_in[239]
  PIN w0_mask_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 333.050 0.800 333.350 ;
    END
  END w0_mask_in[240]
  PIN w0_mask_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 334.410 0.800 334.710 ;
    END
  END w0_mask_in[241]
  PIN w0_mask_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 335.770 0.800 336.070 ;
    END
  END w0_mask_in[242]
  PIN w0_mask_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 337.130 0.800 337.430 ;
    END
  END w0_mask_in[243]
  PIN w0_mask_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 338.490 0.800 338.790 ;
    END
  END w0_mask_in[244]
  PIN w0_mask_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 339.850 0.800 340.150 ;
    END
  END w0_mask_in[245]
  PIN w0_mask_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 341.210 0.800 341.510 ;
    END
  END w0_mask_in[246]
  PIN w0_mask_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 342.570 0.800 342.870 ;
    END
  END w0_mask_in[247]
  PIN w0_mask_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 343.930 0.800 344.230 ;
    END
  END w0_mask_in[248]
  PIN w0_mask_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 345.290 0.800 345.590 ;
    END
  END w0_mask_in[249]
  PIN w0_mask_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 346.650 0.800 346.950 ;
    END
  END w0_mask_in[250]
  PIN w0_mask_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 348.010 0.800 348.310 ;
    END
  END w0_mask_in[251]
  PIN w0_mask_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 349.370 0.800 349.670 ;
    END
  END w0_mask_in[252]
  PIN w0_mask_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 350.730 0.800 351.030 ;
    END
  END w0_mask_in[253]
  PIN w0_mask_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 352.090 0.800 352.390 ;
    END
  END w0_mask_in[254]
  PIN w0_mask_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 353.450 0.800 353.750 ;
    END
  END w0_mask_in[255]
  PIN w0_mask_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 354.810 0.800 355.110 ;
    END
  END w0_mask_in[256]
  PIN w0_mask_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 356.170 0.800 356.470 ;
    END
  END w0_mask_in[257]
  PIN w0_mask_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 357.530 0.800 357.830 ;
    END
  END w0_mask_in[258]
  PIN w0_mask_in[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 358.890 0.800 359.190 ;
    END
  END w0_mask_in[259]
  PIN w0_mask_in[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 360.250 0.800 360.550 ;
    END
  END w0_mask_in[260]
  PIN w0_mask_in[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 361.610 0.800 361.910 ;
    END
  END w0_mask_in[261]
  PIN w0_mask_in[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 362.970 0.800 363.270 ;
    END
  END w0_mask_in[262]
  PIN w0_mask_in[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 364.330 0.800 364.630 ;
    END
  END w0_mask_in[263]
  PIN w0_mask_in[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 365.690 0.800 365.990 ;
    END
  END w0_mask_in[264]
  PIN w0_mask_in[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 367.050 0.800 367.350 ;
    END
  END w0_mask_in[265]
  PIN w0_mask_in[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 368.410 0.800 368.710 ;
    END
  END w0_mask_in[266]
  PIN w0_mask_in[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 369.770 0.800 370.070 ;
    END
  END w0_mask_in[267]
  PIN w0_mask_in[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 371.130 0.800 371.430 ;
    END
  END w0_mask_in[268]
  PIN w0_mask_in[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 372.490 0.800 372.790 ;
    END
  END w0_mask_in[269]
  PIN w0_mask_in[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 373.850 0.800 374.150 ;
    END
  END w0_mask_in[270]
  PIN w0_mask_in[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 375.210 0.800 375.510 ;
    END
  END w0_mask_in[271]
  PIN w0_mask_in[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 376.570 0.800 376.870 ;
    END
  END w0_mask_in[272]
  PIN w0_mask_in[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 377.930 0.800 378.230 ;
    END
  END w0_mask_in[273]
  PIN w0_mask_in[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 379.290 0.800 379.590 ;
    END
  END w0_mask_in[274]
  PIN w0_mask_in[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 380.650 0.800 380.950 ;
    END
  END w0_mask_in[275]
  PIN w0_mask_in[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 382.010 0.800 382.310 ;
    END
  END w0_mask_in[276]
  PIN w0_mask_in[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 383.370 0.800 383.670 ;
    END
  END w0_mask_in[277]
  PIN w0_mask_in[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 384.730 0.800 385.030 ;
    END
  END w0_mask_in[278]
  PIN w0_mask_in[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 386.090 0.800 386.390 ;
    END
  END w0_mask_in[279]
  PIN w0_mask_in[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 387.450 0.800 387.750 ;
    END
  END w0_mask_in[280]
  PIN w0_mask_in[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 388.810 0.800 389.110 ;
    END
  END w0_mask_in[281]
  PIN w0_mask_in[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 390.170 0.800 390.470 ;
    END
  END w0_mask_in[282]
  PIN w0_mask_in[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 391.530 0.800 391.830 ;
    END
  END w0_mask_in[283]
  PIN w0_mask_in[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 392.890 0.800 393.190 ;
    END
  END w0_mask_in[284]
  PIN w0_mask_in[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 394.250 0.800 394.550 ;
    END
  END w0_mask_in[285]
  PIN w0_mask_in[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 395.610 0.800 395.910 ;
    END
  END w0_mask_in[286]
  PIN w0_mask_in[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 396.970 0.800 397.270 ;
    END
  END w0_mask_in[287]
  PIN w0_mask_in[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 398.330 0.800 398.630 ;
    END
  END w0_mask_in[288]
  PIN w0_mask_in[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 399.690 0.800 399.990 ;
    END
  END w0_mask_in[289]
  PIN w0_mask_in[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 401.050 0.800 401.350 ;
    END
  END w0_mask_in[290]
  PIN w0_mask_in[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 402.410 0.800 402.710 ;
    END
  END w0_mask_in[291]
  PIN w0_mask_in[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 403.770 0.800 404.070 ;
    END
  END w0_mask_in[292]
  PIN w0_mask_in[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 405.130 0.800 405.430 ;
    END
  END w0_mask_in[293]
  PIN w0_mask_in[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 406.490 0.800 406.790 ;
    END
  END w0_mask_in[294]
  PIN w0_mask_in[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 407.850 0.800 408.150 ;
    END
  END w0_mask_in[295]
  PIN w0_mask_in[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 409.210 0.800 409.510 ;
    END
  END w0_mask_in[296]
  PIN w0_mask_in[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 410.570 0.800 410.870 ;
    END
  END w0_mask_in[297]
  PIN w0_mask_in[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 411.930 0.800 412.230 ;
    END
  END w0_mask_in[298]
  PIN w0_mask_in[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 413.290 0.800 413.590 ;
    END
  END w0_mask_in[299]
  PIN w0_mask_in[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 414.650 0.800 414.950 ;
    END
  END w0_mask_in[300]
  PIN w0_mask_in[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 416.010 0.800 416.310 ;
    END
  END w0_mask_in[301]
  PIN w0_mask_in[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 417.370 0.800 417.670 ;
    END
  END w0_mask_in[302]
  PIN w0_mask_in[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 418.730 0.800 419.030 ;
    END
  END w0_mask_in[303]
  PIN w0_mask_in[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 420.090 0.800 420.390 ;
    END
  END w0_mask_in[304]
  PIN w0_mask_in[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 421.450 0.800 421.750 ;
    END
  END w0_mask_in[305]
  PIN w0_mask_in[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 422.810 0.800 423.110 ;
    END
  END w0_mask_in[306]
  PIN w0_mask_in[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 424.170 0.800 424.470 ;
    END
  END w0_mask_in[307]
  PIN w0_mask_in[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 425.530 0.800 425.830 ;
    END
  END w0_mask_in[308]
  PIN w0_mask_in[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 426.890 0.800 427.190 ;
    END
  END w0_mask_in[309]
  PIN w0_mask_in[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 428.250 0.800 428.550 ;
    END
  END w0_mask_in[310]
  PIN w0_mask_in[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 429.610 0.800 429.910 ;
    END
  END w0_mask_in[311]
  PIN w0_mask_in[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 430.970 0.800 431.270 ;
    END
  END w0_mask_in[312]
  PIN w0_mask_in[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 432.330 0.800 432.630 ;
    END
  END w0_mask_in[313]
  PIN w0_mask_in[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 433.690 0.800 433.990 ;
    END
  END w0_mask_in[314]
  PIN w0_mask_in[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 435.050 0.800 435.350 ;
    END
  END w0_mask_in[315]
  PIN w0_mask_in[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 436.410 0.800 436.710 ;
    END
  END w0_mask_in[316]
  PIN w0_mask_in[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 437.770 0.800 438.070 ;
    END
  END w0_mask_in[317]
  PIN w0_mask_in[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 439.130 0.800 439.430 ;
    END
  END w0_mask_in[318]
  PIN w0_mask_in[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 440.490 0.800 440.790 ;
    END
  END w0_mask_in[319]
  PIN w0_mask_in[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 441.850 0.800 442.150 ;
    END
  END w0_mask_in[320]
  PIN w0_mask_in[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 443.210 0.800 443.510 ;
    END
  END w0_mask_in[321]
  PIN w0_mask_in[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 444.570 0.800 444.870 ;
    END
  END w0_mask_in[322]
  PIN w0_mask_in[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 445.930 0.800 446.230 ;
    END
  END w0_mask_in[323]
  PIN w0_mask_in[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 447.290 0.800 447.590 ;
    END
  END w0_mask_in[324]
  PIN w0_mask_in[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 448.650 0.800 448.950 ;
    END
  END w0_mask_in[325]
  PIN w0_mask_in[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 450.010 0.800 450.310 ;
    END
  END w0_mask_in[326]
  PIN w0_mask_in[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 451.370 0.800 451.670 ;
    END
  END w0_mask_in[327]
  PIN w0_mask_in[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 452.730 0.800 453.030 ;
    END
  END w0_mask_in[328]
  PIN w0_mask_in[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 454.090 0.800 454.390 ;
    END
  END w0_mask_in[329]
  PIN w0_mask_in[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 455.450 0.800 455.750 ;
    END
  END w0_mask_in[330]
  PIN w0_mask_in[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 456.810 0.800 457.110 ;
    END
  END w0_mask_in[331]
  PIN w0_mask_in[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 458.170 0.800 458.470 ;
    END
  END w0_mask_in[332]
  PIN w0_mask_in[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 459.530 0.800 459.830 ;
    END
  END w0_mask_in[333]
  PIN w0_mask_in[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 460.890 0.800 461.190 ;
    END
  END w0_mask_in[334]
  PIN w0_mask_in[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 462.250 0.800 462.550 ;
    END
  END w0_mask_in[335]
  PIN w0_mask_in[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 463.610 0.800 463.910 ;
    END
  END w0_mask_in[336]
  PIN w0_mask_in[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 464.970 0.800 465.270 ;
    END
  END w0_mask_in[337]
  PIN w0_mask_in[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 466.330 0.800 466.630 ;
    END
  END w0_mask_in[338]
  PIN w0_mask_in[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 467.690 0.800 467.990 ;
    END
  END w0_mask_in[339]
  PIN w0_mask_in[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 469.050 0.800 469.350 ;
    END
  END w0_mask_in[340]
  PIN w0_mask_in[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 470.410 0.800 470.710 ;
    END
  END w0_mask_in[341]
  PIN w0_mask_in[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 471.770 0.800 472.070 ;
    END
  END w0_mask_in[342]
  PIN w0_mask_in[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 473.130 0.800 473.430 ;
    END
  END w0_mask_in[343]
  PIN w0_mask_in[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 474.490 0.800 474.790 ;
    END
  END w0_mask_in[344]
  PIN w0_mask_in[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 475.850 0.800 476.150 ;
    END
  END w0_mask_in[345]
  PIN w0_mask_in[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 477.210 0.800 477.510 ;
    END
  END w0_mask_in[346]
  PIN w0_mask_in[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 478.570 0.800 478.870 ;
    END
  END w0_mask_in[347]
  PIN w0_mask_in[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 479.930 0.800 480.230 ;
    END
  END w0_mask_in[348]
  PIN w0_mask_in[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 481.290 0.800 481.590 ;
    END
  END w0_mask_in[349]
  PIN w0_mask_in[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 482.650 0.800 482.950 ;
    END
  END w0_mask_in[350]
  PIN w0_mask_in[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 484.010 0.800 484.310 ;
    END
  END w0_mask_in[351]
  PIN w0_mask_in[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 485.370 0.800 485.670 ;
    END
  END w0_mask_in[352]
  PIN w0_mask_in[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 486.730 0.800 487.030 ;
    END
  END w0_mask_in[353]
  PIN w0_mask_in[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 488.090 0.800 488.390 ;
    END
  END w0_mask_in[354]
  PIN w0_mask_in[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 489.450 0.800 489.750 ;
    END
  END w0_mask_in[355]
  PIN w0_mask_in[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 490.810 0.800 491.110 ;
    END
  END w0_mask_in[356]
  PIN w0_mask_in[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 492.170 0.800 492.470 ;
    END
  END w0_mask_in[357]
  PIN w0_mask_in[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 493.530 0.800 493.830 ;
    END
  END w0_mask_in[358]
  PIN w0_mask_in[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 494.890 0.800 495.190 ;
    END
  END w0_mask_in[359]
  PIN w0_mask_in[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 496.250 0.800 496.550 ;
    END
  END w0_mask_in[360]
  PIN w0_mask_in[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 497.610 0.800 497.910 ;
    END
  END w0_mask_in[361]
  PIN w0_mask_in[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 498.970 0.800 499.270 ;
    END
  END w0_mask_in[362]
  PIN w0_mask_in[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 500.330 0.800 500.630 ;
    END
  END w0_mask_in[363]
  PIN w0_mask_in[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 501.690 0.800 501.990 ;
    END
  END w0_mask_in[364]
  PIN w0_mask_in[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 503.050 0.800 503.350 ;
    END
  END w0_mask_in[365]
  PIN w0_mask_in[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 504.410 0.800 504.710 ;
    END
  END w0_mask_in[366]
  PIN w0_mask_in[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 505.770 0.800 506.070 ;
    END
  END w0_mask_in[367]
  PIN w0_mask_in[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 507.130 0.800 507.430 ;
    END
  END w0_mask_in[368]
  PIN w0_mask_in[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 508.490 0.800 508.790 ;
    END
  END w0_mask_in[369]
  PIN w0_mask_in[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 509.850 0.800 510.150 ;
    END
  END w0_mask_in[370]
  PIN w0_mask_in[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 511.210 0.800 511.510 ;
    END
  END w0_mask_in[371]
  PIN w0_mask_in[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 512.570 0.800 512.870 ;
    END
  END w0_mask_in[372]
  PIN w0_mask_in[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 513.930 0.800 514.230 ;
    END
  END w0_mask_in[373]
  PIN w0_mask_in[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 515.290 0.800 515.590 ;
    END
  END w0_mask_in[374]
  PIN w0_mask_in[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 516.650 0.800 516.950 ;
    END
  END w0_mask_in[375]
  PIN w0_mask_in[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 518.010 0.800 518.310 ;
    END
  END w0_mask_in[376]
  PIN w0_mask_in[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 519.370 0.800 519.670 ;
    END
  END w0_mask_in[377]
  PIN w0_mask_in[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 520.730 0.800 521.030 ;
    END
  END w0_mask_in[378]
  PIN w0_mask_in[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 522.090 0.800 522.390 ;
    END
  END w0_mask_in[379]
  PIN w0_mask_in[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 523.450 0.800 523.750 ;
    END
  END w0_mask_in[380]
  PIN w0_mask_in[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 524.810 0.800 525.110 ;
    END
  END w0_mask_in[381]
  PIN w0_mask_in[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 526.170 0.800 526.470 ;
    END
  END w0_mask_in[382]
  PIN w0_mask_in[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 527.530 0.800 527.830 ;
    END
  END w0_mask_in[383]
  PIN w0_mask_in[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 528.890 0.800 529.190 ;
    END
  END w0_mask_in[384]
  PIN w0_mask_in[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 530.250 0.800 530.550 ;
    END
  END w0_mask_in[385]
  PIN w0_mask_in[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 531.610 0.800 531.910 ;
    END
  END w0_mask_in[386]
  PIN w0_mask_in[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 532.970 0.800 533.270 ;
    END
  END w0_mask_in[387]
  PIN w0_mask_in[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 534.330 0.800 534.630 ;
    END
  END w0_mask_in[388]
  PIN w0_mask_in[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 535.690 0.800 535.990 ;
    END
  END w0_mask_in[389]
  PIN w0_mask_in[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 537.050 0.800 537.350 ;
    END
  END w0_mask_in[390]
  PIN w0_mask_in[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 538.410 0.800 538.710 ;
    END
  END w0_mask_in[391]
  PIN w0_mask_in[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 539.770 0.800 540.070 ;
    END
  END w0_mask_in[392]
  PIN w0_mask_in[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 541.130 0.800 541.430 ;
    END
  END w0_mask_in[393]
  PIN w0_mask_in[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 542.490 0.800 542.790 ;
    END
  END w0_mask_in[394]
  PIN w0_mask_in[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 543.850 0.800 544.150 ;
    END
  END w0_mask_in[395]
  PIN w0_mask_in[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 545.210 0.800 545.510 ;
    END
  END w0_mask_in[396]
  PIN w0_mask_in[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 546.570 0.800 546.870 ;
    END
  END w0_mask_in[397]
  PIN w0_mask_in[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 547.930 0.800 548.230 ;
    END
  END w0_mask_in[398]
  PIN w0_mask_in[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 549.290 0.800 549.590 ;
    END
  END w0_mask_in[399]
  PIN w0_mask_in[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 550.650 0.800 550.950 ;
    END
  END w0_mask_in[400]
  PIN w0_mask_in[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 552.010 0.800 552.310 ;
    END
  END w0_mask_in[401]
  PIN w0_mask_in[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 553.370 0.800 553.670 ;
    END
  END w0_mask_in[402]
  PIN w0_mask_in[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 554.730 0.800 555.030 ;
    END
  END w0_mask_in[403]
  PIN w0_mask_in[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 556.090 0.800 556.390 ;
    END
  END w0_mask_in[404]
  PIN w0_mask_in[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 557.450 0.800 557.750 ;
    END
  END w0_mask_in[405]
  PIN w0_mask_in[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 558.810 0.800 559.110 ;
    END
  END w0_mask_in[406]
  PIN w0_mask_in[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 560.170 0.800 560.470 ;
    END
  END w0_mask_in[407]
  PIN w0_mask_in[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 561.530 0.800 561.830 ;
    END
  END w0_mask_in[408]
  PIN w0_mask_in[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 562.890 0.800 563.190 ;
    END
  END w0_mask_in[409]
  PIN w0_mask_in[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 564.250 0.800 564.550 ;
    END
  END w0_mask_in[410]
  PIN w0_mask_in[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 565.610 0.800 565.910 ;
    END
  END w0_mask_in[411]
  PIN w0_mask_in[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 566.970 0.800 567.270 ;
    END
  END w0_mask_in[412]
  PIN w0_mask_in[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 568.330 0.800 568.630 ;
    END
  END w0_mask_in[413]
  PIN w0_mask_in[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 569.690 0.800 569.990 ;
    END
  END w0_mask_in[414]
  PIN w0_mask_in[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 571.050 0.800 571.350 ;
    END
  END w0_mask_in[415]
  PIN w0_mask_in[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 572.410 0.800 572.710 ;
    END
  END w0_mask_in[416]
  PIN w0_mask_in[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 573.770 0.800 574.070 ;
    END
  END w0_mask_in[417]
  PIN w0_mask_in[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 575.130 0.800 575.430 ;
    END
  END w0_mask_in[418]
  PIN w0_mask_in[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 576.490 0.800 576.790 ;
    END
  END w0_mask_in[419]
  PIN w0_mask_in[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 577.850 0.800 578.150 ;
    END
  END w0_mask_in[420]
  PIN w0_mask_in[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 579.210 0.800 579.510 ;
    END
  END w0_mask_in[421]
  PIN w0_mask_in[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 580.570 0.800 580.870 ;
    END
  END w0_mask_in[422]
  PIN w0_mask_in[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 581.930 0.800 582.230 ;
    END
  END w0_mask_in[423]
  PIN w0_mask_in[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 583.290 0.800 583.590 ;
    END
  END w0_mask_in[424]
  PIN w0_mask_in[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 584.650 0.800 584.950 ;
    END
  END w0_mask_in[425]
  PIN w0_mask_in[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 586.010 0.800 586.310 ;
    END
  END w0_mask_in[426]
  PIN w0_mask_in[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 587.370 0.800 587.670 ;
    END
  END w0_mask_in[427]
  PIN w0_mask_in[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 588.730 0.800 589.030 ;
    END
  END w0_mask_in[428]
  PIN w0_mask_in[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 590.090 0.800 590.390 ;
    END
  END w0_mask_in[429]
  PIN w0_mask_in[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 591.450 0.800 591.750 ;
    END
  END w0_mask_in[430]
  PIN w0_mask_in[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 592.810 0.800 593.110 ;
    END
  END w0_mask_in[431]
  PIN w0_mask_in[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 594.170 0.800 594.470 ;
    END
  END w0_mask_in[432]
  PIN w0_mask_in[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 595.530 0.800 595.830 ;
    END
  END w0_mask_in[433]
  PIN w0_mask_in[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 596.890 0.800 597.190 ;
    END
  END w0_mask_in[434]
  PIN w0_mask_in[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 598.250 0.800 598.550 ;
    END
  END w0_mask_in[435]
  PIN w0_mask_in[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 599.610 0.800 599.910 ;
    END
  END w0_mask_in[436]
  PIN w0_mask_in[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 600.970 0.800 601.270 ;
    END
  END w0_mask_in[437]
  PIN w0_mask_in[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 602.330 0.800 602.630 ;
    END
  END w0_mask_in[438]
  PIN w0_mask_in[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 603.690 0.800 603.990 ;
    END
  END w0_mask_in[439]
  PIN w0_mask_in[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 605.050 0.800 605.350 ;
    END
  END w0_mask_in[440]
  PIN w0_mask_in[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 606.410 0.800 606.710 ;
    END
  END w0_mask_in[441]
  PIN w0_mask_in[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 607.770 0.800 608.070 ;
    END
  END w0_mask_in[442]
  PIN w0_mask_in[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 609.130 0.800 609.430 ;
    END
  END w0_mask_in[443]
  PIN w0_mask_in[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 610.490 0.800 610.790 ;
    END
  END w0_mask_in[444]
  PIN w0_mask_in[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 611.850 0.800 612.150 ;
    END
  END w0_mask_in[445]
  PIN w0_mask_in[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 613.210 0.800 613.510 ;
    END
  END w0_mask_in[446]
  PIN w0_mask_in[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 614.570 0.800 614.870 ;
    END
  END w0_mask_in[447]
  PIN w0_mask_in[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 615.930 0.800 616.230 ;
    END
  END w0_mask_in[448]
  PIN w0_mask_in[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 617.290 0.800 617.590 ;
    END
  END w0_mask_in[449]
  PIN w0_mask_in[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 618.650 0.800 618.950 ;
    END
  END w0_mask_in[450]
  PIN w0_mask_in[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 620.010 0.800 620.310 ;
    END
  END w0_mask_in[451]
  PIN w0_mask_in[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 621.370 0.800 621.670 ;
    END
  END w0_mask_in[452]
  PIN w0_mask_in[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 622.730 0.800 623.030 ;
    END
  END w0_mask_in[453]
  PIN w0_mask_in[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 624.090 0.800 624.390 ;
    END
  END w0_mask_in[454]
  PIN w0_mask_in[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 625.450 0.800 625.750 ;
    END
  END w0_mask_in[455]
  PIN w0_mask_in[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 626.810 0.800 627.110 ;
    END
  END w0_mask_in[456]
  PIN w0_mask_in[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 628.170 0.800 628.470 ;
    END
  END w0_mask_in[457]
  PIN w0_mask_in[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 629.530 0.800 629.830 ;
    END
  END w0_mask_in[458]
  PIN w0_mask_in[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 630.890 0.800 631.190 ;
    END
  END w0_mask_in[459]
  PIN w0_mask_in[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 632.250 0.800 632.550 ;
    END
  END w0_mask_in[460]
  PIN w0_mask_in[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 633.610 0.800 633.910 ;
    END
  END w0_mask_in[461]
  PIN w0_mask_in[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 634.970 0.800 635.270 ;
    END
  END w0_mask_in[462]
  PIN w0_mask_in[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 636.330 0.800 636.630 ;
    END
  END w0_mask_in[463]
  PIN w0_mask_in[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 637.690 0.800 637.990 ;
    END
  END w0_mask_in[464]
  PIN w0_mask_in[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 639.050 0.800 639.350 ;
    END
  END w0_mask_in[465]
  PIN w0_mask_in[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 640.410 0.800 640.710 ;
    END
  END w0_mask_in[466]
  PIN w0_mask_in[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 641.770 0.800 642.070 ;
    END
  END w0_mask_in[467]
  PIN w0_mask_in[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 643.130 0.800 643.430 ;
    END
  END w0_mask_in[468]
  PIN w0_mask_in[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 644.490 0.800 644.790 ;
    END
  END w0_mask_in[469]
  PIN w0_mask_in[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 645.850 0.800 646.150 ;
    END
  END w0_mask_in[470]
  PIN w0_mask_in[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 647.210 0.800 647.510 ;
    END
  END w0_mask_in[471]
  PIN w0_mask_in[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 648.570 0.800 648.870 ;
    END
  END w0_mask_in[472]
  PIN w0_mask_in[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 649.930 0.800 650.230 ;
    END
  END w0_mask_in[473]
  PIN w0_mask_in[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 651.290 0.800 651.590 ;
    END
  END w0_mask_in[474]
  PIN w0_mask_in[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 652.650 0.800 652.950 ;
    END
  END w0_mask_in[475]
  PIN w0_mask_in[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 654.010 0.800 654.310 ;
    END
  END w0_mask_in[476]
  PIN w0_mask_in[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 655.370 0.800 655.670 ;
    END
  END w0_mask_in[477]
  PIN w0_mask_in[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 656.730 0.800 657.030 ;
    END
  END w0_mask_in[478]
  PIN w0_mask_in[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 658.090 0.800 658.390 ;
    END
  END w0_mask_in[479]
  PIN w0_mask_in[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 659.450 0.800 659.750 ;
    END
  END w0_mask_in[480]
  PIN w0_mask_in[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 660.810 0.800 661.110 ;
    END
  END w0_mask_in[481]
  PIN w0_mask_in[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 662.170 0.800 662.470 ;
    END
  END w0_mask_in[482]
  PIN w0_mask_in[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 663.530 0.800 663.830 ;
    END
  END w0_mask_in[483]
  PIN w0_mask_in[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 664.890 0.800 665.190 ;
    END
  END w0_mask_in[484]
  PIN w0_mask_in[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 666.250 0.800 666.550 ;
    END
  END w0_mask_in[485]
  PIN w0_mask_in[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 667.610 0.800 667.910 ;
    END
  END w0_mask_in[486]
  PIN w0_mask_in[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 668.970 0.800 669.270 ;
    END
  END w0_mask_in[487]
  PIN w0_mask_in[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 670.330 0.800 670.630 ;
    END
  END w0_mask_in[488]
  PIN w0_mask_in[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 671.690 0.800 671.990 ;
    END
  END w0_mask_in[489]
  PIN w0_mask_in[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 673.050 0.800 673.350 ;
    END
  END w0_mask_in[490]
  PIN w0_mask_in[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 674.410 0.800 674.710 ;
    END
  END w0_mask_in[491]
  PIN w0_mask_in[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 675.770 0.800 676.070 ;
    END
  END w0_mask_in[492]
  PIN w0_mask_in[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 677.130 0.800 677.430 ;
    END
  END w0_mask_in[493]
  PIN w0_mask_in[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 678.490 0.800 678.790 ;
    END
  END w0_mask_in[494]
  PIN w0_mask_in[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 679.850 0.800 680.150 ;
    END
  END w0_mask_in[495]
  PIN w0_mask_in[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 681.210 0.800 681.510 ;
    END
  END w0_mask_in[496]
  PIN w0_mask_in[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 682.570 0.800 682.870 ;
    END
  END w0_mask_in[497]
  PIN w0_mask_in[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 683.930 0.800 684.230 ;
    END
  END w0_mask_in[498]
  PIN w0_mask_in[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 685.290 0.800 685.590 ;
    END
  END w0_mask_in[499]
  PIN w0_mask_in[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 686.650 0.800 686.950 ;
    END
  END w0_mask_in[500]
  PIN w0_mask_in[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 688.010 0.800 688.310 ;
    END
  END w0_mask_in[501]
  PIN w0_mask_in[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 689.370 0.800 689.670 ;
    END
  END w0_mask_in[502]
  PIN w0_mask_in[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 690.730 0.800 691.030 ;
    END
  END w0_mask_in[503]
  PIN w0_mask_in[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 692.090 0.800 692.390 ;
    END
  END w0_mask_in[504]
  PIN w0_mask_in[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 693.450 0.800 693.750 ;
    END
  END w0_mask_in[505]
  PIN w0_mask_in[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 694.810 0.800 695.110 ;
    END
  END w0_mask_in[506]
  PIN w0_mask_in[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 696.170 0.800 696.470 ;
    END
  END w0_mask_in[507]
  PIN w0_mask_in[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 697.530 0.800 697.830 ;
    END
  END w0_mask_in[508]
  PIN w0_mask_in[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 698.890 0.800 699.190 ;
    END
  END w0_mask_in[509]
  PIN w0_mask_in[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 700.250 0.800 700.550 ;
    END
  END w0_mask_in[510]
  PIN w0_mask_in[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 701.610 0.800 701.910 ;
    END
  END w0_mask_in[511]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 783.210 0.800 783.510 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 784.570 0.800 784.870 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 785.930 0.800 786.230 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 787.290 0.800 787.590 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 788.650 0.800 788.950 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 790.010 0.800 790.310 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 791.370 0.800 791.670 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 792.730 0.800 793.030 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 794.090 0.800 794.390 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 795.450 0.800 795.750 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 796.810 0.800 797.110 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 798.170 0.800 798.470 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 799.530 0.800 799.830 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 800.890 0.800 801.190 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 802.250 0.800 802.550 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 803.610 0.800 803.910 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 804.970 0.800 805.270 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 806.330 0.800 806.630 ;
    END
  END w0_wd_in[17]
  PIN w0_wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 807.690 0.800 807.990 ;
    END
  END w0_wd_in[18]
  PIN w0_wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 809.050 0.800 809.350 ;
    END
  END w0_wd_in[19]
  PIN w0_wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 810.410 0.800 810.710 ;
    END
  END w0_wd_in[20]
  PIN w0_wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 811.770 0.800 812.070 ;
    END
  END w0_wd_in[21]
  PIN w0_wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 813.130 0.800 813.430 ;
    END
  END w0_wd_in[22]
  PIN w0_wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 814.490 0.800 814.790 ;
    END
  END w0_wd_in[23]
  PIN w0_wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 815.850 0.800 816.150 ;
    END
  END w0_wd_in[24]
  PIN w0_wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 817.210 0.800 817.510 ;
    END
  END w0_wd_in[25]
  PIN w0_wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 818.570 0.800 818.870 ;
    END
  END w0_wd_in[26]
  PIN w0_wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 819.930 0.800 820.230 ;
    END
  END w0_wd_in[27]
  PIN w0_wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 821.290 0.800 821.590 ;
    END
  END w0_wd_in[28]
  PIN w0_wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 822.650 0.800 822.950 ;
    END
  END w0_wd_in[29]
  PIN w0_wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 824.010 0.800 824.310 ;
    END
  END w0_wd_in[30]
  PIN w0_wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 825.370 0.800 825.670 ;
    END
  END w0_wd_in[31]
  PIN w0_wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 826.730 0.800 827.030 ;
    END
  END w0_wd_in[32]
  PIN w0_wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 828.090 0.800 828.390 ;
    END
  END w0_wd_in[33]
  PIN w0_wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 829.450 0.800 829.750 ;
    END
  END w0_wd_in[34]
  PIN w0_wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 830.810 0.800 831.110 ;
    END
  END w0_wd_in[35]
  PIN w0_wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 832.170 0.800 832.470 ;
    END
  END w0_wd_in[36]
  PIN w0_wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 833.530 0.800 833.830 ;
    END
  END w0_wd_in[37]
  PIN w0_wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 834.890 0.800 835.190 ;
    END
  END w0_wd_in[38]
  PIN w0_wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 836.250 0.800 836.550 ;
    END
  END w0_wd_in[39]
  PIN w0_wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 837.610 0.800 837.910 ;
    END
  END w0_wd_in[40]
  PIN w0_wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 838.970 0.800 839.270 ;
    END
  END w0_wd_in[41]
  PIN w0_wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 840.330 0.800 840.630 ;
    END
  END w0_wd_in[42]
  PIN w0_wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 841.690 0.800 841.990 ;
    END
  END w0_wd_in[43]
  PIN w0_wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 843.050 0.800 843.350 ;
    END
  END w0_wd_in[44]
  PIN w0_wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 844.410 0.800 844.710 ;
    END
  END w0_wd_in[45]
  PIN w0_wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 845.770 0.800 846.070 ;
    END
  END w0_wd_in[46]
  PIN w0_wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 847.130 0.800 847.430 ;
    END
  END w0_wd_in[47]
  PIN w0_wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 848.490 0.800 848.790 ;
    END
  END w0_wd_in[48]
  PIN w0_wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 849.850 0.800 850.150 ;
    END
  END w0_wd_in[49]
  PIN w0_wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 851.210 0.800 851.510 ;
    END
  END w0_wd_in[50]
  PIN w0_wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 852.570 0.800 852.870 ;
    END
  END w0_wd_in[51]
  PIN w0_wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 853.930 0.800 854.230 ;
    END
  END w0_wd_in[52]
  PIN w0_wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 855.290 0.800 855.590 ;
    END
  END w0_wd_in[53]
  PIN w0_wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 856.650 0.800 856.950 ;
    END
  END w0_wd_in[54]
  PIN w0_wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 858.010 0.800 858.310 ;
    END
  END w0_wd_in[55]
  PIN w0_wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 859.370 0.800 859.670 ;
    END
  END w0_wd_in[56]
  PIN w0_wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 860.730 0.800 861.030 ;
    END
  END w0_wd_in[57]
  PIN w0_wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 862.090 0.800 862.390 ;
    END
  END w0_wd_in[58]
  PIN w0_wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 863.450 0.800 863.750 ;
    END
  END w0_wd_in[59]
  PIN w0_wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 864.810 0.800 865.110 ;
    END
  END w0_wd_in[60]
  PIN w0_wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 866.170 0.800 866.470 ;
    END
  END w0_wd_in[61]
  PIN w0_wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 867.530 0.800 867.830 ;
    END
  END w0_wd_in[62]
  PIN w0_wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 868.890 0.800 869.190 ;
    END
  END w0_wd_in[63]
  PIN w0_wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 870.250 0.800 870.550 ;
    END
  END w0_wd_in[64]
  PIN w0_wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 871.610 0.800 871.910 ;
    END
  END w0_wd_in[65]
  PIN w0_wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 872.970 0.800 873.270 ;
    END
  END w0_wd_in[66]
  PIN w0_wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 874.330 0.800 874.630 ;
    END
  END w0_wd_in[67]
  PIN w0_wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 875.690 0.800 875.990 ;
    END
  END w0_wd_in[68]
  PIN w0_wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 877.050 0.800 877.350 ;
    END
  END w0_wd_in[69]
  PIN w0_wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 878.410 0.800 878.710 ;
    END
  END w0_wd_in[70]
  PIN w0_wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 879.770 0.800 880.070 ;
    END
  END w0_wd_in[71]
  PIN w0_wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 881.130 0.800 881.430 ;
    END
  END w0_wd_in[72]
  PIN w0_wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 882.490 0.800 882.790 ;
    END
  END w0_wd_in[73]
  PIN w0_wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 883.850 0.800 884.150 ;
    END
  END w0_wd_in[74]
  PIN w0_wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 885.210 0.800 885.510 ;
    END
  END w0_wd_in[75]
  PIN w0_wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 886.570 0.800 886.870 ;
    END
  END w0_wd_in[76]
  PIN w0_wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 887.930 0.800 888.230 ;
    END
  END w0_wd_in[77]
  PIN w0_wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 889.290 0.800 889.590 ;
    END
  END w0_wd_in[78]
  PIN w0_wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 890.650 0.800 890.950 ;
    END
  END w0_wd_in[79]
  PIN w0_wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 892.010 0.800 892.310 ;
    END
  END w0_wd_in[80]
  PIN w0_wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 893.370 0.800 893.670 ;
    END
  END w0_wd_in[81]
  PIN w0_wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 894.730 0.800 895.030 ;
    END
  END w0_wd_in[82]
  PIN w0_wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 896.090 0.800 896.390 ;
    END
  END w0_wd_in[83]
  PIN w0_wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 897.450 0.800 897.750 ;
    END
  END w0_wd_in[84]
  PIN w0_wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 898.810 0.800 899.110 ;
    END
  END w0_wd_in[85]
  PIN w0_wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 900.170 0.800 900.470 ;
    END
  END w0_wd_in[86]
  PIN w0_wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 901.530 0.800 901.830 ;
    END
  END w0_wd_in[87]
  PIN w0_wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 902.890 0.800 903.190 ;
    END
  END w0_wd_in[88]
  PIN w0_wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 904.250 0.800 904.550 ;
    END
  END w0_wd_in[89]
  PIN w0_wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 905.610 0.800 905.910 ;
    END
  END w0_wd_in[90]
  PIN w0_wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 906.970 0.800 907.270 ;
    END
  END w0_wd_in[91]
  PIN w0_wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 908.330 0.800 908.630 ;
    END
  END w0_wd_in[92]
  PIN w0_wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 909.690 0.800 909.990 ;
    END
  END w0_wd_in[93]
  PIN w0_wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 911.050 0.800 911.350 ;
    END
  END w0_wd_in[94]
  PIN w0_wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 912.410 0.800 912.710 ;
    END
  END w0_wd_in[95]
  PIN w0_wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 913.770 0.800 914.070 ;
    END
  END w0_wd_in[96]
  PIN w0_wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 915.130 0.800 915.430 ;
    END
  END w0_wd_in[97]
  PIN w0_wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 916.490 0.800 916.790 ;
    END
  END w0_wd_in[98]
  PIN w0_wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 917.850 0.800 918.150 ;
    END
  END w0_wd_in[99]
  PIN w0_wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 919.210 0.800 919.510 ;
    END
  END w0_wd_in[100]
  PIN w0_wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 920.570 0.800 920.870 ;
    END
  END w0_wd_in[101]
  PIN w0_wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 921.930 0.800 922.230 ;
    END
  END w0_wd_in[102]
  PIN w0_wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 923.290 0.800 923.590 ;
    END
  END w0_wd_in[103]
  PIN w0_wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 924.650 0.800 924.950 ;
    END
  END w0_wd_in[104]
  PIN w0_wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 926.010 0.800 926.310 ;
    END
  END w0_wd_in[105]
  PIN w0_wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 927.370 0.800 927.670 ;
    END
  END w0_wd_in[106]
  PIN w0_wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 928.730 0.800 929.030 ;
    END
  END w0_wd_in[107]
  PIN w0_wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 930.090 0.800 930.390 ;
    END
  END w0_wd_in[108]
  PIN w0_wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 931.450 0.800 931.750 ;
    END
  END w0_wd_in[109]
  PIN w0_wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 932.810 0.800 933.110 ;
    END
  END w0_wd_in[110]
  PIN w0_wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 934.170 0.800 934.470 ;
    END
  END w0_wd_in[111]
  PIN w0_wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 935.530 0.800 935.830 ;
    END
  END w0_wd_in[112]
  PIN w0_wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 936.890 0.800 937.190 ;
    END
  END w0_wd_in[113]
  PIN w0_wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 938.250 0.800 938.550 ;
    END
  END w0_wd_in[114]
  PIN w0_wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 939.610 0.800 939.910 ;
    END
  END w0_wd_in[115]
  PIN w0_wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 940.970 0.800 941.270 ;
    END
  END w0_wd_in[116]
  PIN w0_wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 942.330 0.800 942.630 ;
    END
  END w0_wd_in[117]
  PIN w0_wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 943.690 0.800 943.990 ;
    END
  END w0_wd_in[118]
  PIN w0_wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 945.050 0.800 945.350 ;
    END
  END w0_wd_in[119]
  PIN w0_wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 946.410 0.800 946.710 ;
    END
  END w0_wd_in[120]
  PIN w0_wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 947.770 0.800 948.070 ;
    END
  END w0_wd_in[121]
  PIN w0_wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 949.130 0.800 949.430 ;
    END
  END w0_wd_in[122]
  PIN w0_wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 950.490 0.800 950.790 ;
    END
  END w0_wd_in[123]
  PIN w0_wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 951.850 0.800 952.150 ;
    END
  END w0_wd_in[124]
  PIN w0_wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 953.210 0.800 953.510 ;
    END
  END w0_wd_in[125]
  PIN w0_wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 954.570 0.800 954.870 ;
    END
  END w0_wd_in[126]
  PIN w0_wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 955.930 0.800 956.230 ;
    END
  END w0_wd_in[127]
  PIN w0_wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 957.290 0.800 957.590 ;
    END
  END w0_wd_in[128]
  PIN w0_wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 958.650 0.800 958.950 ;
    END
  END w0_wd_in[129]
  PIN w0_wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 960.010 0.800 960.310 ;
    END
  END w0_wd_in[130]
  PIN w0_wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 961.370 0.800 961.670 ;
    END
  END w0_wd_in[131]
  PIN w0_wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 962.730 0.800 963.030 ;
    END
  END w0_wd_in[132]
  PIN w0_wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 964.090 0.800 964.390 ;
    END
  END w0_wd_in[133]
  PIN w0_wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 965.450 0.800 965.750 ;
    END
  END w0_wd_in[134]
  PIN w0_wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 966.810 0.800 967.110 ;
    END
  END w0_wd_in[135]
  PIN w0_wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 968.170 0.800 968.470 ;
    END
  END w0_wd_in[136]
  PIN w0_wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 969.530 0.800 969.830 ;
    END
  END w0_wd_in[137]
  PIN w0_wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 970.890 0.800 971.190 ;
    END
  END w0_wd_in[138]
  PIN w0_wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 972.250 0.800 972.550 ;
    END
  END w0_wd_in[139]
  PIN w0_wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 973.610 0.800 973.910 ;
    END
  END w0_wd_in[140]
  PIN w0_wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 974.970 0.800 975.270 ;
    END
  END w0_wd_in[141]
  PIN w0_wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 976.330 0.800 976.630 ;
    END
  END w0_wd_in[142]
  PIN w0_wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 977.690 0.800 977.990 ;
    END
  END w0_wd_in[143]
  PIN w0_wd_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 979.050 0.800 979.350 ;
    END
  END w0_wd_in[144]
  PIN w0_wd_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 980.410 0.800 980.710 ;
    END
  END w0_wd_in[145]
  PIN w0_wd_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 981.770 0.800 982.070 ;
    END
  END w0_wd_in[146]
  PIN w0_wd_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 983.130 0.800 983.430 ;
    END
  END w0_wd_in[147]
  PIN w0_wd_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 984.490 0.800 984.790 ;
    END
  END w0_wd_in[148]
  PIN w0_wd_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 985.850 0.800 986.150 ;
    END
  END w0_wd_in[149]
  PIN w0_wd_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 987.210 0.800 987.510 ;
    END
  END w0_wd_in[150]
  PIN w0_wd_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 988.570 0.800 988.870 ;
    END
  END w0_wd_in[151]
  PIN w0_wd_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 989.930 0.800 990.230 ;
    END
  END w0_wd_in[152]
  PIN w0_wd_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 991.290 0.800 991.590 ;
    END
  END w0_wd_in[153]
  PIN w0_wd_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 992.650 0.800 992.950 ;
    END
  END w0_wd_in[154]
  PIN w0_wd_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 994.010 0.800 994.310 ;
    END
  END w0_wd_in[155]
  PIN w0_wd_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 995.370 0.800 995.670 ;
    END
  END w0_wd_in[156]
  PIN w0_wd_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 996.730 0.800 997.030 ;
    END
  END w0_wd_in[157]
  PIN w0_wd_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 998.090 0.800 998.390 ;
    END
  END w0_wd_in[158]
  PIN w0_wd_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 999.450 0.800 999.750 ;
    END
  END w0_wd_in[159]
  PIN w0_wd_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1000.810 0.800 1001.110 ;
    END
  END w0_wd_in[160]
  PIN w0_wd_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1002.170 0.800 1002.470 ;
    END
  END w0_wd_in[161]
  PIN w0_wd_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1003.530 0.800 1003.830 ;
    END
  END w0_wd_in[162]
  PIN w0_wd_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1004.890 0.800 1005.190 ;
    END
  END w0_wd_in[163]
  PIN w0_wd_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1006.250 0.800 1006.550 ;
    END
  END w0_wd_in[164]
  PIN w0_wd_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1007.610 0.800 1007.910 ;
    END
  END w0_wd_in[165]
  PIN w0_wd_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1008.970 0.800 1009.270 ;
    END
  END w0_wd_in[166]
  PIN w0_wd_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1010.330 0.800 1010.630 ;
    END
  END w0_wd_in[167]
  PIN w0_wd_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1011.690 0.800 1011.990 ;
    END
  END w0_wd_in[168]
  PIN w0_wd_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1013.050 0.800 1013.350 ;
    END
  END w0_wd_in[169]
  PIN w0_wd_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1014.410 0.800 1014.710 ;
    END
  END w0_wd_in[170]
  PIN w0_wd_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1015.770 0.800 1016.070 ;
    END
  END w0_wd_in[171]
  PIN w0_wd_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1017.130 0.800 1017.430 ;
    END
  END w0_wd_in[172]
  PIN w0_wd_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1018.490 0.800 1018.790 ;
    END
  END w0_wd_in[173]
  PIN w0_wd_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1019.850 0.800 1020.150 ;
    END
  END w0_wd_in[174]
  PIN w0_wd_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1021.210 0.800 1021.510 ;
    END
  END w0_wd_in[175]
  PIN w0_wd_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1022.570 0.800 1022.870 ;
    END
  END w0_wd_in[176]
  PIN w0_wd_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1023.930 0.800 1024.230 ;
    END
  END w0_wd_in[177]
  PIN w0_wd_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1025.290 0.800 1025.590 ;
    END
  END w0_wd_in[178]
  PIN w0_wd_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1026.650 0.800 1026.950 ;
    END
  END w0_wd_in[179]
  PIN w0_wd_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1028.010 0.800 1028.310 ;
    END
  END w0_wd_in[180]
  PIN w0_wd_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1029.370 0.800 1029.670 ;
    END
  END w0_wd_in[181]
  PIN w0_wd_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1030.730 0.800 1031.030 ;
    END
  END w0_wd_in[182]
  PIN w0_wd_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1032.090 0.800 1032.390 ;
    END
  END w0_wd_in[183]
  PIN w0_wd_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1033.450 0.800 1033.750 ;
    END
  END w0_wd_in[184]
  PIN w0_wd_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1034.810 0.800 1035.110 ;
    END
  END w0_wd_in[185]
  PIN w0_wd_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1036.170 0.800 1036.470 ;
    END
  END w0_wd_in[186]
  PIN w0_wd_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1037.530 0.800 1037.830 ;
    END
  END w0_wd_in[187]
  PIN w0_wd_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1038.890 0.800 1039.190 ;
    END
  END w0_wd_in[188]
  PIN w0_wd_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1040.250 0.800 1040.550 ;
    END
  END w0_wd_in[189]
  PIN w0_wd_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1041.610 0.800 1041.910 ;
    END
  END w0_wd_in[190]
  PIN w0_wd_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1042.970 0.800 1043.270 ;
    END
  END w0_wd_in[191]
  PIN w0_wd_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1044.330 0.800 1044.630 ;
    END
  END w0_wd_in[192]
  PIN w0_wd_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1045.690 0.800 1045.990 ;
    END
  END w0_wd_in[193]
  PIN w0_wd_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1047.050 0.800 1047.350 ;
    END
  END w0_wd_in[194]
  PIN w0_wd_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1048.410 0.800 1048.710 ;
    END
  END w0_wd_in[195]
  PIN w0_wd_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1049.770 0.800 1050.070 ;
    END
  END w0_wd_in[196]
  PIN w0_wd_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1051.130 0.800 1051.430 ;
    END
  END w0_wd_in[197]
  PIN w0_wd_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1052.490 0.800 1052.790 ;
    END
  END w0_wd_in[198]
  PIN w0_wd_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1053.850 0.800 1054.150 ;
    END
  END w0_wd_in[199]
  PIN w0_wd_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1055.210 0.800 1055.510 ;
    END
  END w0_wd_in[200]
  PIN w0_wd_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1056.570 0.800 1056.870 ;
    END
  END w0_wd_in[201]
  PIN w0_wd_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1057.930 0.800 1058.230 ;
    END
  END w0_wd_in[202]
  PIN w0_wd_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1059.290 0.800 1059.590 ;
    END
  END w0_wd_in[203]
  PIN w0_wd_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1060.650 0.800 1060.950 ;
    END
  END w0_wd_in[204]
  PIN w0_wd_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1062.010 0.800 1062.310 ;
    END
  END w0_wd_in[205]
  PIN w0_wd_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1063.370 0.800 1063.670 ;
    END
  END w0_wd_in[206]
  PIN w0_wd_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1064.730 0.800 1065.030 ;
    END
  END w0_wd_in[207]
  PIN w0_wd_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1066.090 0.800 1066.390 ;
    END
  END w0_wd_in[208]
  PIN w0_wd_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1067.450 0.800 1067.750 ;
    END
  END w0_wd_in[209]
  PIN w0_wd_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1068.810 0.800 1069.110 ;
    END
  END w0_wd_in[210]
  PIN w0_wd_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1070.170 0.800 1070.470 ;
    END
  END w0_wd_in[211]
  PIN w0_wd_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1071.530 0.800 1071.830 ;
    END
  END w0_wd_in[212]
  PIN w0_wd_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1072.890 0.800 1073.190 ;
    END
  END w0_wd_in[213]
  PIN w0_wd_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1074.250 0.800 1074.550 ;
    END
  END w0_wd_in[214]
  PIN w0_wd_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1075.610 0.800 1075.910 ;
    END
  END w0_wd_in[215]
  PIN w0_wd_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1076.970 0.800 1077.270 ;
    END
  END w0_wd_in[216]
  PIN w0_wd_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1078.330 0.800 1078.630 ;
    END
  END w0_wd_in[217]
  PIN w0_wd_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1079.690 0.800 1079.990 ;
    END
  END w0_wd_in[218]
  PIN w0_wd_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1081.050 0.800 1081.350 ;
    END
  END w0_wd_in[219]
  PIN w0_wd_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1082.410 0.800 1082.710 ;
    END
  END w0_wd_in[220]
  PIN w0_wd_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1083.770 0.800 1084.070 ;
    END
  END w0_wd_in[221]
  PIN w0_wd_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1085.130 0.800 1085.430 ;
    END
  END w0_wd_in[222]
  PIN w0_wd_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1086.490 0.800 1086.790 ;
    END
  END w0_wd_in[223]
  PIN w0_wd_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1087.850 0.800 1088.150 ;
    END
  END w0_wd_in[224]
  PIN w0_wd_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1089.210 0.800 1089.510 ;
    END
  END w0_wd_in[225]
  PIN w0_wd_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1090.570 0.800 1090.870 ;
    END
  END w0_wd_in[226]
  PIN w0_wd_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1091.930 0.800 1092.230 ;
    END
  END w0_wd_in[227]
  PIN w0_wd_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1093.290 0.800 1093.590 ;
    END
  END w0_wd_in[228]
  PIN w0_wd_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1094.650 0.800 1094.950 ;
    END
  END w0_wd_in[229]
  PIN w0_wd_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1096.010 0.800 1096.310 ;
    END
  END w0_wd_in[230]
  PIN w0_wd_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1097.370 0.800 1097.670 ;
    END
  END w0_wd_in[231]
  PIN w0_wd_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1098.730 0.800 1099.030 ;
    END
  END w0_wd_in[232]
  PIN w0_wd_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1100.090 0.800 1100.390 ;
    END
  END w0_wd_in[233]
  PIN w0_wd_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1101.450 0.800 1101.750 ;
    END
  END w0_wd_in[234]
  PIN w0_wd_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1102.810 0.800 1103.110 ;
    END
  END w0_wd_in[235]
  PIN w0_wd_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1104.170 0.800 1104.470 ;
    END
  END w0_wd_in[236]
  PIN w0_wd_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1105.530 0.800 1105.830 ;
    END
  END w0_wd_in[237]
  PIN w0_wd_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1106.890 0.800 1107.190 ;
    END
  END w0_wd_in[238]
  PIN w0_wd_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1108.250 0.800 1108.550 ;
    END
  END w0_wd_in[239]
  PIN w0_wd_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1109.610 0.800 1109.910 ;
    END
  END w0_wd_in[240]
  PIN w0_wd_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1110.970 0.800 1111.270 ;
    END
  END w0_wd_in[241]
  PIN w0_wd_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1112.330 0.800 1112.630 ;
    END
  END w0_wd_in[242]
  PIN w0_wd_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1113.690 0.800 1113.990 ;
    END
  END w0_wd_in[243]
  PIN w0_wd_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1115.050 0.800 1115.350 ;
    END
  END w0_wd_in[244]
  PIN w0_wd_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1116.410 0.800 1116.710 ;
    END
  END w0_wd_in[245]
  PIN w0_wd_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1117.770 0.800 1118.070 ;
    END
  END w0_wd_in[246]
  PIN w0_wd_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1119.130 0.800 1119.430 ;
    END
  END w0_wd_in[247]
  PIN w0_wd_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1120.490 0.800 1120.790 ;
    END
  END w0_wd_in[248]
  PIN w0_wd_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1121.850 0.800 1122.150 ;
    END
  END w0_wd_in[249]
  PIN w0_wd_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1123.210 0.800 1123.510 ;
    END
  END w0_wd_in[250]
  PIN w0_wd_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1124.570 0.800 1124.870 ;
    END
  END w0_wd_in[251]
  PIN w0_wd_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1125.930 0.800 1126.230 ;
    END
  END w0_wd_in[252]
  PIN w0_wd_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1127.290 0.800 1127.590 ;
    END
  END w0_wd_in[253]
  PIN w0_wd_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1128.650 0.800 1128.950 ;
    END
  END w0_wd_in[254]
  PIN w0_wd_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1130.010 0.800 1130.310 ;
    END
  END w0_wd_in[255]
  PIN w0_wd_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1131.370 0.800 1131.670 ;
    END
  END w0_wd_in[256]
  PIN w0_wd_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1132.730 0.800 1133.030 ;
    END
  END w0_wd_in[257]
  PIN w0_wd_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1134.090 0.800 1134.390 ;
    END
  END w0_wd_in[258]
  PIN w0_wd_in[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1135.450 0.800 1135.750 ;
    END
  END w0_wd_in[259]
  PIN w0_wd_in[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1136.810 0.800 1137.110 ;
    END
  END w0_wd_in[260]
  PIN w0_wd_in[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1138.170 0.800 1138.470 ;
    END
  END w0_wd_in[261]
  PIN w0_wd_in[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1139.530 0.800 1139.830 ;
    END
  END w0_wd_in[262]
  PIN w0_wd_in[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1140.890 0.800 1141.190 ;
    END
  END w0_wd_in[263]
  PIN w0_wd_in[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1142.250 0.800 1142.550 ;
    END
  END w0_wd_in[264]
  PIN w0_wd_in[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1143.610 0.800 1143.910 ;
    END
  END w0_wd_in[265]
  PIN w0_wd_in[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1144.970 0.800 1145.270 ;
    END
  END w0_wd_in[266]
  PIN w0_wd_in[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1146.330 0.800 1146.630 ;
    END
  END w0_wd_in[267]
  PIN w0_wd_in[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1147.690 0.800 1147.990 ;
    END
  END w0_wd_in[268]
  PIN w0_wd_in[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1149.050 0.800 1149.350 ;
    END
  END w0_wd_in[269]
  PIN w0_wd_in[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1150.410 0.800 1150.710 ;
    END
  END w0_wd_in[270]
  PIN w0_wd_in[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1151.770 0.800 1152.070 ;
    END
  END w0_wd_in[271]
  PIN w0_wd_in[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1153.130 0.800 1153.430 ;
    END
  END w0_wd_in[272]
  PIN w0_wd_in[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1154.490 0.800 1154.790 ;
    END
  END w0_wd_in[273]
  PIN w0_wd_in[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1155.850 0.800 1156.150 ;
    END
  END w0_wd_in[274]
  PIN w0_wd_in[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1157.210 0.800 1157.510 ;
    END
  END w0_wd_in[275]
  PIN w0_wd_in[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1158.570 0.800 1158.870 ;
    END
  END w0_wd_in[276]
  PIN w0_wd_in[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1159.930 0.800 1160.230 ;
    END
  END w0_wd_in[277]
  PIN w0_wd_in[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1161.290 0.800 1161.590 ;
    END
  END w0_wd_in[278]
  PIN w0_wd_in[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1162.650 0.800 1162.950 ;
    END
  END w0_wd_in[279]
  PIN w0_wd_in[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1164.010 0.800 1164.310 ;
    END
  END w0_wd_in[280]
  PIN w0_wd_in[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1165.370 0.800 1165.670 ;
    END
  END w0_wd_in[281]
  PIN w0_wd_in[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1166.730 0.800 1167.030 ;
    END
  END w0_wd_in[282]
  PIN w0_wd_in[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1168.090 0.800 1168.390 ;
    END
  END w0_wd_in[283]
  PIN w0_wd_in[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1169.450 0.800 1169.750 ;
    END
  END w0_wd_in[284]
  PIN w0_wd_in[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1170.810 0.800 1171.110 ;
    END
  END w0_wd_in[285]
  PIN w0_wd_in[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1172.170 0.800 1172.470 ;
    END
  END w0_wd_in[286]
  PIN w0_wd_in[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1173.530 0.800 1173.830 ;
    END
  END w0_wd_in[287]
  PIN w0_wd_in[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1174.890 0.800 1175.190 ;
    END
  END w0_wd_in[288]
  PIN w0_wd_in[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1176.250 0.800 1176.550 ;
    END
  END w0_wd_in[289]
  PIN w0_wd_in[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1177.610 0.800 1177.910 ;
    END
  END w0_wd_in[290]
  PIN w0_wd_in[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1178.970 0.800 1179.270 ;
    END
  END w0_wd_in[291]
  PIN w0_wd_in[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1180.330 0.800 1180.630 ;
    END
  END w0_wd_in[292]
  PIN w0_wd_in[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1181.690 0.800 1181.990 ;
    END
  END w0_wd_in[293]
  PIN w0_wd_in[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1183.050 0.800 1183.350 ;
    END
  END w0_wd_in[294]
  PIN w0_wd_in[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1184.410 0.800 1184.710 ;
    END
  END w0_wd_in[295]
  PIN w0_wd_in[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1185.770 0.800 1186.070 ;
    END
  END w0_wd_in[296]
  PIN w0_wd_in[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1187.130 0.800 1187.430 ;
    END
  END w0_wd_in[297]
  PIN w0_wd_in[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1188.490 0.800 1188.790 ;
    END
  END w0_wd_in[298]
  PIN w0_wd_in[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1189.850 0.800 1190.150 ;
    END
  END w0_wd_in[299]
  PIN w0_wd_in[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1191.210 0.800 1191.510 ;
    END
  END w0_wd_in[300]
  PIN w0_wd_in[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1192.570 0.800 1192.870 ;
    END
  END w0_wd_in[301]
  PIN w0_wd_in[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1193.930 0.800 1194.230 ;
    END
  END w0_wd_in[302]
  PIN w0_wd_in[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1195.290 0.800 1195.590 ;
    END
  END w0_wd_in[303]
  PIN w0_wd_in[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1196.650 0.800 1196.950 ;
    END
  END w0_wd_in[304]
  PIN w0_wd_in[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1198.010 0.800 1198.310 ;
    END
  END w0_wd_in[305]
  PIN w0_wd_in[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1199.370 0.800 1199.670 ;
    END
  END w0_wd_in[306]
  PIN w0_wd_in[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1200.730 0.800 1201.030 ;
    END
  END w0_wd_in[307]
  PIN w0_wd_in[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1202.090 0.800 1202.390 ;
    END
  END w0_wd_in[308]
  PIN w0_wd_in[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1203.450 0.800 1203.750 ;
    END
  END w0_wd_in[309]
  PIN w0_wd_in[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1204.810 0.800 1205.110 ;
    END
  END w0_wd_in[310]
  PIN w0_wd_in[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1206.170 0.800 1206.470 ;
    END
  END w0_wd_in[311]
  PIN w0_wd_in[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1207.530 0.800 1207.830 ;
    END
  END w0_wd_in[312]
  PIN w0_wd_in[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1208.890 0.800 1209.190 ;
    END
  END w0_wd_in[313]
  PIN w0_wd_in[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1210.250 0.800 1210.550 ;
    END
  END w0_wd_in[314]
  PIN w0_wd_in[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1211.610 0.800 1211.910 ;
    END
  END w0_wd_in[315]
  PIN w0_wd_in[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1212.970 0.800 1213.270 ;
    END
  END w0_wd_in[316]
  PIN w0_wd_in[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1214.330 0.800 1214.630 ;
    END
  END w0_wd_in[317]
  PIN w0_wd_in[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1215.690 0.800 1215.990 ;
    END
  END w0_wd_in[318]
  PIN w0_wd_in[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1217.050 0.800 1217.350 ;
    END
  END w0_wd_in[319]
  PIN w0_wd_in[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1218.410 0.800 1218.710 ;
    END
  END w0_wd_in[320]
  PIN w0_wd_in[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1219.770 0.800 1220.070 ;
    END
  END w0_wd_in[321]
  PIN w0_wd_in[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1221.130 0.800 1221.430 ;
    END
  END w0_wd_in[322]
  PIN w0_wd_in[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1222.490 0.800 1222.790 ;
    END
  END w0_wd_in[323]
  PIN w0_wd_in[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1223.850 0.800 1224.150 ;
    END
  END w0_wd_in[324]
  PIN w0_wd_in[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1225.210 0.800 1225.510 ;
    END
  END w0_wd_in[325]
  PIN w0_wd_in[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1226.570 0.800 1226.870 ;
    END
  END w0_wd_in[326]
  PIN w0_wd_in[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1227.930 0.800 1228.230 ;
    END
  END w0_wd_in[327]
  PIN w0_wd_in[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1229.290 0.800 1229.590 ;
    END
  END w0_wd_in[328]
  PIN w0_wd_in[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1230.650 0.800 1230.950 ;
    END
  END w0_wd_in[329]
  PIN w0_wd_in[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1232.010 0.800 1232.310 ;
    END
  END w0_wd_in[330]
  PIN w0_wd_in[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1233.370 0.800 1233.670 ;
    END
  END w0_wd_in[331]
  PIN w0_wd_in[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1234.730 0.800 1235.030 ;
    END
  END w0_wd_in[332]
  PIN w0_wd_in[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1236.090 0.800 1236.390 ;
    END
  END w0_wd_in[333]
  PIN w0_wd_in[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1237.450 0.800 1237.750 ;
    END
  END w0_wd_in[334]
  PIN w0_wd_in[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1238.810 0.800 1239.110 ;
    END
  END w0_wd_in[335]
  PIN w0_wd_in[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1240.170 0.800 1240.470 ;
    END
  END w0_wd_in[336]
  PIN w0_wd_in[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1241.530 0.800 1241.830 ;
    END
  END w0_wd_in[337]
  PIN w0_wd_in[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1242.890 0.800 1243.190 ;
    END
  END w0_wd_in[338]
  PIN w0_wd_in[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1244.250 0.800 1244.550 ;
    END
  END w0_wd_in[339]
  PIN w0_wd_in[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1245.610 0.800 1245.910 ;
    END
  END w0_wd_in[340]
  PIN w0_wd_in[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1246.970 0.800 1247.270 ;
    END
  END w0_wd_in[341]
  PIN w0_wd_in[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1248.330 0.800 1248.630 ;
    END
  END w0_wd_in[342]
  PIN w0_wd_in[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1249.690 0.800 1249.990 ;
    END
  END w0_wd_in[343]
  PIN w0_wd_in[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1251.050 0.800 1251.350 ;
    END
  END w0_wd_in[344]
  PIN w0_wd_in[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1252.410 0.800 1252.710 ;
    END
  END w0_wd_in[345]
  PIN w0_wd_in[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1253.770 0.800 1254.070 ;
    END
  END w0_wd_in[346]
  PIN w0_wd_in[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1255.130 0.800 1255.430 ;
    END
  END w0_wd_in[347]
  PIN w0_wd_in[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1256.490 0.800 1256.790 ;
    END
  END w0_wd_in[348]
  PIN w0_wd_in[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1257.850 0.800 1258.150 ;
    END
  END w0_wd_in[349]
  PIN w0_wd_in[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1259.210 0.800 1259.510 ;
    END
  END w0_wd_in[350]
  PIN w0_wd_in[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1260.570 0.800 1260.870 ;
    END
  END w0_wd_in[351]
  PIN w0_wd_in[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1261.930 0.800 1262.230 ;
    END
  END w0_wd_in[352]
  PIN w0_wd_in[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1263.290 0.800 1263.590 ;
    END
  END w0_wd_in[353]
  PIN w0_wd_in[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1264.650 0.800 1264.950 ;
    END
  END w0_wd_in[354]
  PIN w0_wd_in[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1266.010 0.800 1266.310 ;
    END
  END w0_wd_in[355]
  PIN w0_wd_in[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1267.370 0.800 1267.670 ;
    END
  END w0_wd_in[356]
  PIN w0_wd_in[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1268.730 0.800 1269.030 ;
    END
  END w0_wd_in[357]
  PIN w0_wd_in[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1270.090 0.800 1270.390 ;
    END
  END w0_wd_in[358]
  PIN w0_wd_in[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1271.450 0.800 1271.750 ;
    END
  END w0_wd_in[359]
  PIN w0_wd_in[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1272.810 0.800 1273.110 ;
    END
  END w0_wd_in[360]
  PIN w0_wd_in[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1274.170 0.800 1274.470 ;
    END
  END w0_wd_in[361]
  PIN w0_wd_in[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1275.530 0.800 1275.830 ;
    END
  END w0_wd_in[362]
  PIN w0_wd_in[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1276.890 0.800 1277.190 ;
    END
  END w0_wd_in[363]
  PIN w0_wd_in[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1278.250 0.800 1278.550 ;
    END
  END w0_wd_in[364]
  PIN w0_wd_in[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1279.610 0.800 1279.910 ;
    END
  END w0_wd_in[365]
  PIN w0_wd_in[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1280.970 0.800 1281.270 ;
    END
  END w0_wd_in[366]
  PIN w0_wd_in[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1282.330 0.800 1282.630 ;
    END
  END w0_wd_in[367]
  PIN w0_wd_in[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1283.690 0.800 1283.990 ;
    END
  END w0_wd_in[368]
  PIN w0_wd_in[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1285.050 0.800 1285.350 ;
    END
  END w0_wd_in[369]
  PIN w0_wd_in[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1286.410 0.800 1286.710 ;
    END
  END w0_wd_in[370]
  PIN w0_wd_in[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1287.770 0.800 1288.070 ;
    END
  END w0_wd_in[371]
  PIN w0_wd_in[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1289.130 0.800 1289.430 ;
    END
  END w0_wd_in[372]
  PIN w0_wd_in[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1290.490 0.800 1290.790 ;
    END
  END w0_wd_in[373]
  PIN w0_wd_in[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1291.850 0.800 1292.150 ;
    END
  END w0_wd_in[374]
  PIN w0_wd_in[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1293.210 0.800 1293.510 ;
    END
  END w0_wd_in[375]
  PIN w0_wd_in[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1294.570 0.800 1294.870 ;
    END
  END w0_wd_in[376]
  PIN w0_wd_in[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1295.930 0.800 1296.230 ;
    END
  END w0_wd_in[377]
  PIN w0_wd_in[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1297.290 0.800 1297.590 ;
    END
  END w0_wd_in[378]
  PIN w0_wd_in[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1298.650 0.800 1298.950 ;
    END
  END w0_wd_in[379]
  PIN w0_wd_in[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1300.010 0.800 1300.310 ;
    END
  END w0_wd_in[380]
  PIN w0_wd_in[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1301.370 0.800 1301.670 ;
    END
  END w0_wd_in[381]
  PIN w0_wd_in[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1302.730 0.800 1303.030 ;
    END
  END w0_wd_in[382]
  PIN w0_wd_in[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1304.090 0.800 1304.390 ;
    END
  END w0_wd_in[383]
  PIN w0_wd_in[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1305.450 0.800 1305.750 ;
    END
  END w0_wd_in[384]
  PIN w0_wd_in[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1306.810 0.800 1307.110 ;
    END
  END w0_wd_in[385]
  PIN w0_wd_in[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1308.170 0.800 1308.470 ;
    END
  END w0_wd_in[386]
  PIN w0_wd_in[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1309.530 0.800 1309.830 ;
    END
  END w0_wd_in[387]
  PIN w0_wd_in[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1310.890 0.800 1311.190 ;
    END
  END w0_wd_in[388]
  PIN w0_wd_in[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1312.250 0.800 1312.550 ;
    END
  END w0_wd_in[389]
  PIN w0_wd_in[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1313.610 0.800 1313.910 ;
    END
  END w0_wd_in[390]
  PIN w0_wd_in[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1314.970 0.800 1315.270 ;
    END
  END w0_wd_in[391]
  PIN w0_wd_in[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1316.330 0.800 1316.630 ;
    END
  END w0_wd_in[392]
  PIN w0_wd_in[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1317.690 0.800 1317.990 ;
    END
  END w0_wd_in[393]
  PIN w0_wd_in[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1319.050 0.800 1319.350 ;
    END
  END w0_wd_in[394]
  PIN w0_wd_in[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1320.410 0.800 1320.710 ;
    END
  END w0_wd_in[395]
  PIN w0_wd_in[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1321.770 0.800 1322.070 ;
    END
  END w0_wd_in[396]
  PIN w0_wd_in[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1323.130 0.800 1323.430 ;
    END
  END w0_wd_in[397]
  PIN w0_wd_in[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1324.490 0.800 1324.790 ;
    END
  END w0_wd_in[398]
  PIN w0_wd_in[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1325.850 0.800 1326.150 ;
    END
  END w0_wd_in[399]
  PIN w0_wd_in[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1327.210 0.800 1327.510 ;
    END
  END w0_wd_in[400]
  PIN w0_wd_in[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1328.570 0.800 1328.870 ;
    END
  END w0_wd_in[401]
  PIN w0_wd_in[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1329.930 0.800 1330.230 ;
    END
  END w0_wd_in[402]
  PIN w0_wd_in[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1331.290 0.800 1331.590 ;
    END
  END w0_wd_in[403]
  PIN w0_wd_in[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1332.650 0.800 1332.950 ;
    END
  END w0_wd_in[404]
  PIN w0_wd_in[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1334.010 0.800 1334.310 ;
    END
  END w0_wd_in[405]
  PIN w0_wd_in[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1335.370 0.800 1335.670 ;
    END
  END w0_wd_in[406]
  PIN w0_wd_in[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1336.730 0.800 1337.030 ;
    END
  END w0_wd_in[407]
  PIN w0_wd_in[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1338.090 0.800 1338.390 ;
    END
  END w0_wd_in[408]
  PIN w0_wd_in[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1339.450 0.800 1339.750 ;
    END
  END w0_wd_in[409]
  PIN w0_wd_in[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1340.810 0.800 1341.110 ;
    END
  END w0_wd_in[410]
  PIN w0_wd_in[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1342.170 0.800 1342.470 ;
    END
  END w0_wd_in[411]
  PIN w0_wd_in[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1343.530 0.800 1343.830 ;
    END
  END w0_wd_in[412]
  PIN w0_wd_in[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1344.890 0.800 1345.190 ;
    END
  END w0_wd_in[413]
  PIN w0_wd_in[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1346.250 0.800 1346.550 ;
    END
  END w0_wd_in[414]
  PIN w0_wd_in[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1347.610 0.800 1347.910 ;
    END
  END w0_wd_in[415]
  PIN w0_wd_in[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1348.970 0.800 1349.270 ;
    END
  END w0_wd_in[416]
  PIN w0_wd_in[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1350.330 0.800 1350.630 ;
    END
  END w0_wd_in[417]
  PIN w0_wd_in[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1351.690 0.800 1351.990 ;
    END
  END w0_wd_in[418]
  PIN w0_wd_in[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1353.050 0.800 1353.350 ;
    END
  END w0_wd_in[419]
  PIN w0_wd_in[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1354.410 0.800 1354.710 ;
    END
  END w0_wd_in[420]
  PIN w0_wd_in[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1355.770 0.800 1356.070 ;
    END
  END w0_wd_in[421]
  PIN w0_wd_in[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1357.130 0.800 1357.430 ;
    END
  END w0_wd_in[422]
  PIN w0_wd_in[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1358.490 0.800 1358.790 ;
    END
  END w0_wd_in[423]
  PIN w0_wd_in[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1359.850 0.800 1360.150 ;
    END
  END w0_wd_in[424]
  PIN w0_wd_in[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1361.210 0.800 1361.510 ;
    END
  END w0_wd_in[425]
  PIN w0_wd_in[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1362.570 0.800 1362.870 ;
    END
  END w0_wd_in[426]
  PIN w0_wd_in[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1363.930 0.800 1364.230 ;
    END
  END w0_wd_in[427]
  PIN w0_wd_in[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1365.290 0.800 1365.590 ;
    END
  END w0_wd_in[428]
  PIN w0_wd_in[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1366.650 0.800 1366.950 ;
    END
  END w0_wd_in[429]
  PIN w0_wd_in[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1368.010 0.800 1368.310 ;
    END
  END w0_wd_in[430]
  PIN w0_wd_in[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1369.370 0.800 1369.670 ;
    END
  END w0_wd_in[431]
  PIN w0_wd_in[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1370.730 0.800 1371.030 ;
    END
  END w0_wd_in[432]
  PIN w0_wd_in[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1372.090 0.800 1372.390 ;
    END
  END w0_wd_in[433]
  PIN w0_wd_in[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1373.450 0.800 1373.750 ;
    END
  END w0_wd_in[434]
  PIN w0_wd_in[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1374.810 0.800 1375.110 ;
    END
  END w0_wd_in[435]
  PIN w0_wd_in[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1376.170 0.800 1376.470 ;
    END
  END w0_wd_in[436]
  PIN w0_wd_in[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1377.530 0.800 1377.830 ;
    END
  END w0_wd_in[437]
  PIN w0_wd_in[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1378.890 0.800 1379.190 ;
    END
  END w0_wd_in[438]
  PIN w0_wd_in[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1380.250 0.800 1380.550 ;
    END
  END w0_wd_in[439]
  PIN w0_wd_in[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1381.610 0.800 1381.910 ;
    END
  END w0_wd_in[440]
  PIN w0_wd_in[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1382.970 0.800 1383.270 ;
    END
  END w0_wd_in[441]
  PIN w0_wd_in[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1384.330 0.800 1384.630 ;
    END
  END w0_wd_in[442]
  PIN w0_wd_in[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1385.690 0.800 1385.990 ;
    END
  END w0_wd_in[443]
  PIN w0_wd_in[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1387.050 0.800 1387.350 ;
    END
  END w0_wd_in[444]
  PIN w0_wd_in[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1388.410 0.800 1388.710 ;
    END
  END w0_wd_in[445]
  PIN w0_wd_in[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1389.770 0.800 1390.070 ;
    END
  END w0_wd_in[446]
  PIN w0_wd_in[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1391.130 0.800 1391.430 ;
    END
  END w0_wd_in[447]
  PIN w0_wd_in[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1392.490 0.800 1392.790 ;
    END
  END w0_wd_in[448]
  PIN w0_wd_in[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1393.850 0.800 1394.150 ;
    END
  END w0_wd_in[449]
  PIN w0_wd_in[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1395.210 0.800 1395.510 ;
    END
  END w0_wd_in[450]
  PIN w0_wd_in[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1396.570 0.800 1396.870 ;
    END
  END w0_wd_in[451]
  PIN w0_wd_in[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1397.930 0.800 1398.230 ;
    END
  END w0_wd_in[452]
  PIN w0_wd_in[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1399.290 0.800 1399.590 ;
    END
  END w0_wd_in[453]
  PIN w0_wd_in[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1400.650 0.800 1400.950 ;
    END
  END w0_wd_in[454]
  PIN w0_wd_in[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1402.010 0.800 1402.310 ;
    END
  END w0_wd_in[455]
  PIN w0_wd_in[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1403.370 0.800 1403.670 ;
    END
  END w0_wd_in[456]
  PIN w0_wd_in[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1404.730 0.800 1405.030 ;
    END
  END w0_wd_in[457]
  PIN w0_wd_in[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1406.090 0.800 1406.390 ;
    END
  END w0_wd_in[458]
  PIN w0_wd_in[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1407.450 0.800 1407.750 ;
    END
  END w0_wd_in[459]
  PIN w0_wd_in[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1408.810 0.800 1409.110 ;
    END
  END w0_wd_in[460]
  PIN w0_wd_in[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1410.170 0.800 1410.470 ;
    END
  END w0_wd_in[461]
  PIN w0_wd_in[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1411.530 0.800 1411.830 ;
    END
  END w0_wd_in[462]
  PIN w0_wd_in[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1412.890 0.800 1413.190 ;
    END
  END w0_wd_in[463]
  PIN w0_wd_in[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1414.250 0.800 1414.550 ;
    END
  END w0_wd_in[464]
  PIN w0_wd_in[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1415.610 0.800 1415.910 ;
    END
  END w0_wd_in[465]
  PIN w0_wd_in[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1416.970 0.800 1417.270 ;
    END
  END w0_wd_in[466]
  PIN w0_wd_in[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1418.330 0.800 1418.630 ;
    END
  END w0_wd_in[467]
  PIN w0_wd_in[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1419.690 0.800 1419.990 ;
    END
  END w0_wd_in[468]
  PIN w0_wd_in[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1421.050 0.800 1421.350 ;
    END
  END w0_wd_in[469]
  PIN w0_wd_in[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1422.410 0.800 1422.710 ;
    END
  END w0_wd_in[470]
  PIN w0_wd_in[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1423.770 0.800 1424.070 ;
    END
  END w0_wd_in[471]
  PIN w0_wd_in[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1425.130 0.800 1425.430 ;
    END
  END w0_wd_in[472]
  PIN w0_wd_in[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1426.490 0.800 1426.790 ;
    END
  END w0_wd_in[473]
  PIN w0_wd_in[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1427.850 0.800 1428.150 ;
    END
  END w0_wd_in[474]
  PIN w0_wd_in[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1429.210 0.800 1429.510 ;
    END
  END w0_wd_in[475]
  PIN w0_wd_in[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1430.570 0.800 1430.870 ;
    END
  END w0_wd_in[476]
  PIN w0_wd_in[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1431.930 0.800 1432.230 ;
    END
  END w0_wd_in[477]
  PIN w0_wd_in[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1433.290 0.800 1433.590 ;
    END
  END w0_wd_in[478]
  PIN w0_wd_in[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1434.650 0.800 1434.950 ;
    END
  END w0_wd_in[479]
  PIN w0_wd_in[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1436.010 0.800 1436.310 ;
    END
  END w0_wd_in[480]
  PIN w0_wd_in[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1437.370 0.800 1437.670 ;
    END
  END w0_wd_in[481]
  PIN w0_wd_in[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1438.730 0.800 1439.030 ;
    END
  END w0_wd_in[482]
  PIN w0_wd_in[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1440.090 0.800 1440.390 ;
    END
  END w0_wd_in[483]
  PIN w0_wd_in[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1441.450 0.800 1441.750 ;
    END
  END w0_wd_in[484]
  PIN w0_wd_in[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1442.810 0.800 1443.110 ;
    END
  END w0_wd_in[485]
  PIN w0_wd_in[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1444.170 0.800 1444.470 ;
    END
  END w0_wd_in[486]
  PIN w0_wd_in[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1445.530 0.800 1445.830 ;
    END
  END w0_wd_in[487]
  PIN w0_wd_in[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1446.890 0.800 1447.190 ;
    END
  END w0_wd_in[488]
  PIN w0_wd_in[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1448.250 0.800 1448.550 ;
    END
  END w0_wd_in[489]
  PIN w0_wd_in[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1449.610 0.800 1449.910 ;
    END
  END w0_wd_in[490]
  PIN w0_wd_in[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1450.970 0.800 1451.270 ;
    END
  END w0_wd_in[491]
  PIN w0_wd_in[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1452.330 0.800 1452.630 ;
    END
  END w0_wd_in[492]
  PIN w0_wd_in[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1453.690 0.800 1453.990 ;
    END
  END w0_wd_in[493]
  PIN w0_wd_in[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1455.050 0.800 1455.350 ;
    END
  END w0_wd_in[494]
  PIN w0_wd_in[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1456.410 0.800 1456.710 ;
    END
  END w0_wd_in[495]
  PIN w0_wd_in[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1457.770 0.800 1458.070 ;
    END
  END w0_wd_in[496]
  PIN w0_wd_in[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1459.130 0.800 1459.430 ;
    END
  END w0_wd_in[497]
  PIN w0_wd_in[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1460.490 0.800 1460.790 ;
    END
  END w0_wd_in[498]
  PIN w0_wd_in[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1461.850 0.800 1462.150 ;
    END
  END w0_wd_in[499]
  PIN w0_wd_in[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1463.210 0.800 1463.510 ;
    END
  END w0_wd_in[500]
  PIN w0_wd_in[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1464.570 0.800 1464.870 ;
    END
  END w0_wd_in[501]
  PIN w0_wd_in[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1465.930 0.800 1466.230 ;
    END
  END w0_wd_in[502]
  PIN w0_wd_in[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1467.290 0.800 1467.590 ;
    END
  END w0_wd_in[503]
  PIN w0_wd_in[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1468.650 0.800 1468.950 ;
    END
  END w0_wd_in[504]
  PIN w0_wd_in[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1470.010 0.800 1470.310 ;
    END
  END w0_wd_in[505]
  PIN w0_wd_in[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1471.370 0.800 1471.670 ;
    END
  END w0_wd_in[506]
  PIN w0_wd_in[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1472.730 0.800 1473.030 ;
    END
  END w0_wd_in[507]
  PIN w0_wd_in[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1474.090 0.800 1474.390 ;
    END
  END w0_wd_in[508]
  PIN w0_wd_in[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1475.450 0.800 1475.750 ;
    END
  END w0_wd_in[509]
  PIN w0_wd_in[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1476.810 0.800 1477.110 ;
    END
  END w0_wd_in[510]
  PIN w0_wd_in[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1478.170 0.800 1478.470 ;
    END
  END w0_wd_in[511]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 0.000 4.670 0.350 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 6.830 0.000 6.970 0.350 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 9.130 0.000 9.270 0.350 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 11.430 0.000 11.570 0.350 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 13.730 0.000 13.870 0.350 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 16.030 0.000 16.170 0.350 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 18.330 0.000 18.470 0.350 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 20.630 0.000 20.770 0.350 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 22.930 0.000 23.070 0.350 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 25.230 0.000 25.370 0.350 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 27.530 0.000 27.670 0.350 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 29.830 0.000 29.970 0.350 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 32.130 0.000 32.270 0.350 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 34.430 0.000 34.570 0.350 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 36.730 0.000 36.870 0.350 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 39.030 0.000 39.170 0.350 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 41.330 0.000 41.470 0.350 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 43.630 0.000 43.770 0.350 ;
    END
  END r0_rd_out[17]
  PIN r0_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 45.930 0.000 46.070 0.350 ;
    END
  END r0_rd_out[18]
  PIN r0_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 48.230 0.000 48.370 0.350 ;
    END
  END r0_rd_out[19]
  PIN r0_rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 50.530 0.000 50.670 0.350 ;
    END
  END r0_rd_out[20]
  PIN r0_rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 52.830 0.000 52.970 0.350 ;
    END
  END r0_rd_out[21]
  PIN r0_rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 55.130 0.000 55.270 0.350 ;
    END
  END r0_rd_out[22]
  PIN r0_rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 57.430 0.000 57.570 0.350 ;
    END
  END r0_rd_out[23]
  PIN r0_rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 59.730 0.000 59.870 0.350 ;
    END
  END r0_rd_out[24]
  PIN r0_rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 62.030 0.000 62.170 0.350 ;
    END
  END r0_rd_out[25]
  PIN r0_rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 64.330 0.000 64.470 0.350 ;
    END
  END r0_rd_out[26]
  PIN r0_rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 66.630 0.000 66.770 0.350 ;
    END
  END r0_rd_out[27]
  PIN r0_rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 68.930 0.000 69.070 0.350 ;
    END
  END r0_rd_out[28]
  PIN r0_rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 71.230 0.000 71.370 0.350 ;
    END
  END r0_rd_out[29]
  PIN r0_rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 73.530 0.000 73.670 0.350 ;
    END
  END r0_rd_out[30]
  PIN r0_rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 75.830 0.000 75.970 0.350 ;
    END
  END r0_rd_out[31]
  PIN r0_rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 78.130 0.000 78.270 0.350 ;
    END
  END r0_rd_out[32]
  PIN r0_rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 80.430 0.000 80.570 0.350 ;
    END
  END r0_rd_out[33]
  PIN r0_rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 82.730 0.000 82.870 0.350 ;
    END
  END r0_rd_out[34]
  PIN r0_rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 85.030 0.000 85.170 0.350 ;
    END
  END r0_rd_out[35]
  PIN r0_rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 87.330 0.000 87.470 0.350 ;
    END
  END r0_rd_out[36]
  PIN r0_rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 89.630 0.000 89.770 0.350 ;
    END
  END r0_rd_out[37]
  PIN r0_rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 91.930 0.000 92.070 0.350 ;
    END
  END r0_rd_out[38]
  PIN r0_rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 94.230 0.000 94.370 0.350 ;
    END
  END r0_rd_out[39]
  PIN r0_rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 96.530 0.000 96.670 0.350 ;
    END
  END r0_rd_out[40]
  PIN r0_rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 98.830 0.000 98.970 0.350 ;
    END
  END r0_rd_out[41]
  PIN r0_rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 101.130 0.000 101.270 0.350 ;
    END
  END r0_rd_out[42]
  PIN r0_rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 103.430 0.000 103.570 0.350 ;
    END
  END r0_rd_out[43]
  PIN r0_rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 105.730 0.000 105.870 0.350 ;
    END
  END r0_rd_out[44]
  PIN r0_rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 108.030 0.000 108.170 0.350 ;
    END
  END r0_rd_out[45]
  PIN r0_rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 110.330 0.000 110.470 0.350 ;
    END
  END r0_rd_out[46]
  PIN r0_rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 112.630 0.000 112.770 0.350 ;
    END
  END r0_rd_out[47]
  PIN r0_rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 114.930 0.000 115.070 0.350 ;
    END
  END r0_rd_out[48]
  PIN r0_rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 117.230 0.000 117.370 0.350 ;
    END
  END r0_rd_out[49]
  PIN r0_rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 119.530 0.000 119.670 0.350 ;
    END
  END r0_rd_out[50]
  PIN r0_rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 121.830 0.000 121.970 0.350 ;
    END
  END r0_rd_out[51]
  PIN r0_rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 124.130 0.000 124.270 0.350 ;
    END
  END r0_rd_out[52]
  PIN r0_rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 126.430 0.000 126.570 0.350 ;
    END
  END r0_rd_out[53]
  PIN r0_rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 128.730 0.000 128.870 0.350 ;
    END
  END r0_rd_out[54]
  PIN r0_rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 131.030 0.000 131.170 0.350 ;
    END
  END r0_rd_out[55]
  PIN r0_rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 133.330 0.000 133.470 0.350 ;
    END
  END r0_rd_out[56]
  PIN r0_rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 135.630 0.000 135.770 0.350 ;
    END
  END r0_rd_out[57]
  PIN r0_rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 137.930 0.000 138.070 0.350 ;
    END
  END r0_rd_out[58]
  PIN r0_rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 140.230 0.000 140.370 0.350 ;
    END
  END r0_rd_out[59]
  PIN r0_rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 142.530 0.000 142.670 0.350 ;
    END
  END r0_rd_out[60]
  PIN r0_rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 144.830 0.000 144.970 0.350 ;
    END
  END r0_rd_out[61]
  PIN r0_rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 147.130 0.000 147.270 0.350 ;
    END
  END r0_rd_out[62]
  PIN r0_rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 149.430 0.000 149.570 0.350 ;
    END
  END r0_rd_out[63]
  PIN r0_rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 151.730 0.000 151.870 0.350 ;
    END
  END r0_rd_out[64]
  PIN r0_rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 154.030 0.000 154.170 0.350 ;
    END
  END r0_rd_out[65]
  PIN r0_rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 156.330 0.000 156.470 0.350 ;
    END
  END r0_rd_out[66]
  PIN r0_rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 158.630 0.000 158.770 0.350 ;
    END
  END r0_rd_out[67]
  PIN r0_rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 160.930 0.000 161.070 0.350 ;
    END
  END r0_rd_out[68]
  PIN r0_rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 163.230 0.000 163.370 0.350 ;
    END
  END r0_rd_out[69]
  PIN r0_rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 165.530 0.000 165.670 0.350 ;
    END
  END r0_rd_out[70]
  PIN r0_rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 167.830 0.000 167.970 0.350 ;
    END
  END r0_rd_out[71]
  PIN r0_rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 170.130 0.000 170.270 0.350 ;
    END
  END r0_rd_out[72]
  PIN r0_rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 172.430 0.000 172.570 0.350 ;
    END
  END r0_rd_out[73]
  PIN r0_rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 174.730 0.000 174.870 0.350 ;
    END
  END r0_rd_out[74]
  PIN r0_rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 177.030 0.000 177.170 0.350 ;
    END
  END r0_rd_out[75]
  PIN r0_rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 179.330 0.000 179.470 0.350 ;
    END
  END r0_rd_out[76]
  PIN r0_rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 181.630 0.000 181.770 0.350 ;
    END
  END r0_rd_out[77]
  PIN r0_rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 183.930 0.000 184.070 0.350 ;
    END
  END r0_rd_out[78]
  PIN r0_rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 186.230 0.000 186.370 0.350 ;
    END
  END r0_rd_out[79]
  PIN r0_rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 188.530 0.000 188.670 0.350 ;
    END
  END r0_rd_out[80]
  PIN r0_rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 190.830 0.000 190.970 0.350 ;
    END
  END r0_rd_out[81]
  PIN r0_rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 193.130 0.000 193.270 0.350 ;
    END
  END r0_rd_out[82]
  PIN r0_rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 195.430 0.000 195.570 0.350 ;
    END
  END r0_rd_out[83]
  PIN r0_rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 197.730 0.000 197.870 0.350 ;
    END
  END r0_rd_out[84]
  PIN r0_rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 200.030 0.000 200.170 0.350 ;
    END
  END r0_rd_out[85]
  PIN r0_rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 202.330 0.000 202.470 0.350 ;
    END
  END r0_rd_out[86]
  PIN r0_rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 204.630 0.000 204.770 0.350 ;
    END
  END r0_rd_out[87]
  PIN r0_rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 206.930 0.000 207.070 0.350 ;
    END
  END r0_rd_out[88]
  PIN r0_rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 209.230 0.000 209.370 0.350 ;
    END
  END r0_rd_out[89]
  PIN r0_rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 211.530 0.000 211.670 0.350 ;
    END
  END r0_rd_out[90]
  PIN r0_rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 213.830 0.000 213.970 0.350 ;
    END
  END r0_rd_out[91]
  PIN r0_rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 216.130 0.000 216.270 0.350 ;
    END
  END r0_rd_out[92]
  PIN r0_rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 218.430 0.000 218.570 0.350 ;
    END
  END r0_rd_out[93]
  PIN r0_rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 220.730 0.000 220.870 0.350 ;
    END
  END r0_rd_out[94]
  PIN r0_rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 223.030 0.000 223.170 0.350 ;
    END
  END r0_rd_out[95]
  PIN r0_rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 225.330 0.000 225.470 0.350 ;
    END
  END r0_rd_out[96]
  PIN r0_rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 227.630 0.000 227.770 0.350 ;
    END
  END r0_rd_out[97]
  PIN r0_rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 229.930 0.000 230.070 0.350 ;
    END
  END r0_rd_out[98]
  PIN r0_rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 232.230 0.000 232.370 0.350 ;
    END
  END r0_rd_out[99]
  PIN r0_rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 234.530 0.000 234.670 0.350 ;
    END
  END r0_rd_out[100]
  PIN r0_rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 236.830 0.000 236.970 0.350 ;
    END
  END r0_rd_out[101]
  PIN r0_rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 239.130 0.000 239.270 0.350 ;
    END
  END r0_rd_out[102]
  PIN r0_rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 241.430 0.000 241.570 0.350 ;
    END
  END r0_rd_out[103]
  PIN r0_rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 243.730 0.000 243.870 0.350 ;
    END
  END r0_rd_out[104]
  PIN r0_rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 246.030 0.000 246.170 0.350 ;
    END
  END r0_rd_out[105]
  PIN r0_rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 248.330 0.000 248.470 0.350 ;
    END
  END r0_rd_out[106]
  PIN r0_rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 250.630 0.000 250.770 0.350 ;
    END
  END r0_rd_out[107]
  PIN r0_rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 252.930 0.000 253.070 0.350 ;
    END
  END r0_rd_out[108]
  PIN r0_rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 255.230 0.000 255.370 0.350 ;
    END
  END r0_rd_out[109]
  PIN r0_rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 257.530 0.000 257.670 0.350 ;
    END
  END r0_rd_out[110]
  PIN r0_rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 259.830 0.000 259.970 0.350 ;
    END
  END r0_rd_out[111]
  PIN r0_rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 262.130 0.000 262.270 0.350 ;
    END
  END r0_rd_out[112]
  PIN r0_rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 264.430 0.000 264.570 0.350 ;
    END
  END r0_rd_out[113]
  PIN r0_rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 266.730 0.000 266.870 0.350 ;
    END
  END r0_rd_out[114]
  PIN r0_rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 269.030 0.000 269.170 0.350 ;
    END
  END r0_rd_out[115]
  PIN r0_rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 271.330 0.000 271.470 0.350 ;
    END
  END r0_rd_out[116]
  PIN r0_rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 273.630 0.000 273.770 0.350 ;
    END
  END r0_rd_out[117]
  PIN r0_rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 275.930 0.000 276.070 0.350 ;
    END
  END r0_rd_out[118]
  PIN r0_rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 278.230 0.000 278.370 0.350 ;
    END
  END r0_rd_out[119]
  PIN r0_rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 280.530 0.000 280.670 0.350 ;
    END
  END r0_rd_out[120]
  PIN r0_rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 282.830 0.000 282.970 0.350 ;
    END
  END r0_rd_out[121]
  PIN r0_rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 285.130 0.000 285.270 0.350 ;
    END
  END r0_rd_out[122]
  PIN r0_rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 287.430 0.000 287.570 0.350 ;
    END
  END r0_rd_out[123]
  PIN r0_rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 289.730 0.000 289.870 0.350 ;
    END
  END r0_rd_out[124]
  PIN r0_rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 292.030 0.000 292.170 0.350 ;
    END
  END r0_rd_out[125]
  PIN r0_rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 294.330 0.000 294.470 0.350 ;
    END
  END r0_rd_out[126]
  PIN r0_rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 296.630 0.000 296.770 0.350 ;
    END
  END r0_rd_out[127]
  PIN r0_rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 298.930 0.000 299.070 0.350 ;
    END
  END r0_rd_out[128]
  PIN r0_rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 301.230 0.000 301.370 0.350 ;
    END
  END r0_rd_out[129]
  PIN r0_rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 303.530 0.000 303.670 0.350 ;
    END
  END r0_rd_out[130]
  PIN r0_rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 305.830 0.000 305.970 0.350 ;
    END
  END r0_rd_out[131]
  PIN r0_rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 308.130 0.000 308.270 0.350 ;
    END
  END r0_rd_out[132]
  PIN r0_rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 310.430 0.000 310.570 0.350 ;
    END
  END r0_rd_out[133]
  PIN r0_rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 312.730 0.000 312.870 0.350 ;
    END
  END r0_rd_out[134]
  PIN r0_rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 315.030 0.000 315.170 0.350 ;
    END
  END r0_rd_out[135]
  PIN r0_rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 317.330 0.000 317.470 0.350 ;
    END
  END r0_rd_out[136]
  PIN r0_rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 319.630 0.000 319.770 0.350 ;
    END
  END r0_rd_out[137]
  PIN r0_rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 321.930 0.000 322.070 0.350 ;
    END
  END r0_rd_out[138]
  PIN r0_rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 324.230 0.000 324.370 0.350 ;
    END
  END r0_rd_out[139]
  PIN r0_rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 326.530 0.000 326.670 0.350 ;
    END
  END r0_rd_out[140]
  PIN r0_rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 328.830 0.000 328.970 0.350 ;
    END
  END r0_rd_out[141]
  PIN r0_rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 331.130 0.000 331.270 0.350 ;
    END
  END r0_rd_out[142]
  PIN r0_rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 333.430 0.000 333.570 0.350 ;
    END
  END r0_rd_out[143]
  PIN r0_rd_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 335.730 0.000 335.870 0.350 ;
    END
  END r0_rd_out[144]
  PIN r0_rd_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 338.030 0.000 338.170 0.350 ;
    END
  END r0_rd_out[145]
  PIN r0_rd_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 340.330 0.000 340.470 0.350 ;
    END
  END r0_rd_out[146]
  PIN r0_rd_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 342.630 0.000 342.770 0.350 ;
    END
  END r0_rd_out[147]
  PIN r0_rd_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 344.930 0.000 345.070 0.350 ;
    END
  END r0_rd_out[148]
  PIN r0_rd_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 347.230 0.000 347.370 0.350 ;
    END
  END r0_rd_out[149]
  PIN r0_rd_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 349.530 0.000 349.670 0.350 ;
    END
  END r0_rd_out[150]
  PIN r0_rd_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 351.830 0.000 351.970 0.350 ;
    END
  END r0_rd_out[151]
  PIN r0_rd_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 354.130 0.000 354.270 0.350 ;
    END
  END r0_rd_out[152]
  PIN r0_rd_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 356.430 0.000 356.570 0.350 ;
    END
  END r0_rd_out[153]
  PIN r0_rd_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 358.730 0.000 358.870 0.350 ;
    END
  END r0_rd_out[154]
  PIN r0_rd_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 361.030 0.000 361.170 0.350 ;
    END
  END r0_rd_out[155]
  PIN r0_rd_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 363.330 0.000 363.470 0.350 ;
    END
  END r0_rd_out[156]
  PIN r0_rd_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 365.630 0.000 365.770 0.350 ;
    END
  END r0_rd_out[157]
  PIN r0_rd_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 367.930 0.000 368.070 0.350 ;
    END
  END r0_rd_out[158]
  PIN r0_rd_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 370.230 0.000 370.370 0.350 ;
    END
  END r0_rd_out[159]
  PIN r0_rd_out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 372.530 0.000 372.670 0.350 ;
    END
  END r0_rd_out[160]
  PIN r0_rd_out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 374.830 0.000 374.970 0.350 ;
    END
  END r0_rd_out[161]
  PIN r0_rd_out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 377.130 0.000 377.270 0.350 ;
    END
  END r0_rd_out[162]
  PIN r0_rd_out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 379.430 0.000 379.570 0.350 ;
    END
  END r0_rd_out[163]
  PIN r0_rd_out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 381.730 0.000 381.870 0.350 ;
    END
  END r0_rd_out[164]
  PIN r0_rd_out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 384.030 0.000 384.170 0.350 ;
    END
  END r0_rd_out[165]
  PIN r0_rd_out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 386.330 0.000 386.470 0.350 ;
    END
  END r0_rd_out[166]
  PIN r0_rd_out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 388.630 0.000 388.770 0.350 ;
    END
  END r0_rd_out[167]
  PIN r0_rd_out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 390.930 0.000 391.070 0.350 ;
    END
  END r0_rd_out[168]
  PIN r0_rd_out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 393.230 0.000 393.370 0.350 ;
    END
  END r0_rd_out[169]
  PIN r0_rd_out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 395.530 0.000 395.670 0.350 ;
    END
  END r0_rd_out[170]
  PIN r0_rd_out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 397.830 0.000 397.970 0.350 ;
    END
  END r0_rd_out[171]
  PIN r0_rd_out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 400.130 0.000 400.270 0.350 ;
    END
  END r0_rd_out[172]
  PIN r0_rd_out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 402.430 0.000 402.570 0.350 ;
    END
  END r0_rd_out[173]
  PIN r0_rd_out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 404.730 0.000 404.870 0.350 ;
    END
  END r0_rd_out[174]
  PIN r0_rd_out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 407.030 0.000 407.170 0.350 ;
    END
  END r0_rd_out[175]
  PIN r0_rd_out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 409.330 0.000 409.470 0.350 ;
    END
  END r0_rd_out[176]
  PIN r0_rd_out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 411.630 0.000 411.770 0.350 ;
    END
  END r0_rd_out[177]
  PIN r0_rd_out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 413.930 0.000 414.070 0.350 ;
    END
  END r0_rd_out[178]
  PIN r0_rd_out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 416.230 0.000 416.370 0.350 ;
    END
  END r0_rd_out[179]
  PIN r0_rd_out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 418.530 0.000 418.670 0.350 ;
    END
  END r0_rd_out[180]
  PIN r0_rd_out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 420.830 0.000 420.970 0.350 ;
    END
  END r0_rd_out[181]
  PIN r0_rd_out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 423.130 0.000 423.270 0.350 ;
    END
  END r0_rd_out[182]
  PIN r0_rd_out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 425.430 0.000 425.570 0.350 ;
    END
  END r0_rd_out[183]
  PIN r0_rd_out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 427.730 0.000 427.870 0.350 ;
    END
  END r0_rd_out[184]
  PIN r0_rd_out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 430.030 0.000 430.170 0.350 ;
    END
  END r0_rd_out[185]
  PIN r0_rd_out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 432.330 0.000 432.470 0.350 ;
    END
  END r0_rd_out[186]
  PIN r0_rd_out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 434.630 0.000 434.770 0.350 ;
    END
  END r0_rd_out[187]
  PIN r0_rd_out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 436.930 0.000 437.070 0.350 ;
    END
  END r0_rd_out[188]
  PIN r0_rd_out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 439.230 0.000 439.370 0.350 ;
    END
  END r0_rd_out[189]
  PIN r0_rd_out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 441.530 0.000 441.670 0.350 ;
    END
  END r0_rd_out[190]
  PIN r0_rd_out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 443.830 0.000 443.970 0.350 ;
    END
  END r0_rd_out[191]
  PIN r0_rd_out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 446.130 0.000 446.270 0.350 ;
    END
  END r0_rd_out[192]
  PIN r0_rd_out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 448.430 0.000 448.570 0.350 ;
    END
  END r0_rd_out[193]
  PIN r0_rd_out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 450.730 0.000 450.870 0.350 ;
    END
  END r0_rd_out[194]
  PIN r0_rd_out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 453.030 0.000 453.170 0.350 ;
    END
  END r0_rd_out[195]
  PIN r0_rd_out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 455.330 0.000 455.470 0.350 ;
    END
  END r0_rd_out[196]
  PIN r0_rd_out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 457.630 0.000 457.770 0.350 ;
    END
  END r0_rd_out[197]
  PIN r0_rd_out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 459.930 0.000 460.070 0.350 ;
    END
  END r0_rd_out[198]
  PIN r0_rd_out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 462.230 0.000 462.370 0.350 ;
    END
  END r0_rd_out[199]
  PIN r0_rd_out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 464.530 0.000 464.670 0.350 ;
    END
  END r0_rd_out[200]
  PIN r0_rd_out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 466.830 0.000 466.970 0.350 ;
    END
  END r0_rd_out[201]
  PIN r0_rd_out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 469.130 0.000 469.270 0.350 ;
    END
  END r0_rd_out[202]
  PIN r0_rd_out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 471.430 0.000 471.570 0.350 ;
    END
  END r0_rd_out[203]
  PIN r0_rd_out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 473.730 0.000 473.870 0.350 ;
    END
  END r0_rd_out[204]
  PIN r0_rd_out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 476.030 0.000 476.170 0.350 ;
    END
  END r0_rd_out[205]
  PIN r0_rd_out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 478.330 0.000 478.470 0.350 ;
    END
  END r0_rd_out[206]
  PIN r0_rd_out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 480.630 0.000 480.770 0.350 ;
    END
  END r0_rd_out[207]
  PIN r0_rd_out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 482.930 0.000 483.070 0.350 ;
    END
  END r0_rd_out[208]
  PIN r0_rd_out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 485.230 0.000 485.370 0.350 ;
    END
  END r0_rd_out[209]
  PIN r0_rd_out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 487.530 0.000 487.670 0.350 ;
    END
  END r0_rd_out[210]
  PIN r0_rd_out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 489.830 0.000 489.970 0.350 ;
    END
  END r0_rd_out[211]
  PIN r0_rd_out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 492.130 0.000 492.270 0.350 ;
    END
  END r0_rd_out[212]
  PIN r0_rd_out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 494.430 0.000 494.570 0.350 ;
    END
  END r0_rd_out[213]
  PIN r0_rd_out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 496.730 0.000 496.870 0.350 ;
    END
  END r0_rd_out[214]
  PIN r0_rd_out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 499.030 0.000 499.170 0.350 ;
    END
  END r0_rd_out[215]
  PIN r0_rd_out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 501.330 0.000 501.470 0.350 ;
    END
  END r0_rd_out[216]
  PIN r0_rd_out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 503.630 0.000 503.770 0.350 ;
    END
  END r0_rd_out[217]
  PIN r0_rd_out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 505.930 0.000 506.070 0.350 ;
    END
  END r0_rd_out[218]
  PIN r0_rd_out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 508.230 0.000 508.370 0.350 ;
    END
  END r0_rd_out[219]
  PIN r0_rd_out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 510.530 0.000 510.670 0.350 ;
    END
  END r0_rd_out[220]
  PIN r0_rd_out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 512.830 0.000 512.970 0.350 ;
    END
  END r0_rd_out[221]
  PIN r0_rd_out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 515.130 0.000 515.270 0.350 ;
    END
  END r0_rd_out[222]
  PIN r0_rd_out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 517.430 0.000 517.570 0.350 ;
    END
  END r0_rd_out[223]
  PIN r0_rd_out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 519.730 0.000 519.870 0.350 ;
    END
  END r0_rd_out[224]
  PIN r0_rd_out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 522.030 0.000 522.170 0.350 ;
    END
  END r0_rd_out[225]
  PIN r0_rd_out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 524.330 0.000 524.470 0.350 ;
    END
  END r0_rd_out[226]
  PIN r0_rd_out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 526.630 0.000 526.770 0.350 ;
    END
  END r0_rd_out[227]
  PIN r0_rd_out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 528.930 0.000 529.070 0.350 ;
    END
  END r0_rd_out[228]
  PIN r0_rd_out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 531.230 0.000 531.370 0.350 ;
    END
  END r0_rd_out[229]
  PIN r0_rd_out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 533.530 0.000 533.670 0.350 ;
    END
  END r0_rd_out[230]
  PIN r0_rd_out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 535.830 0.000 535.970 0.350 ;
    END
  END r0_rd_out[231]
  PIN r0_rd_out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 538.130 0.000 538.270 0.350 ;
    END
  END r0_rd_out[232]
  PIN r0_rd_out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 540.430 0.000 540.570 0.350 ;
    END
  END r0_rd_out[233]
  PIN r0_rd_out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 542.730 0.000 542.870 0.350 ;
    END
  END r0_rd_out[234]
  PIN r0_rd_out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 545.030 0.000 545.170 0.350 ;
    END
  END r0_rd_out[235]
  PIN r0_rd_out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 547.330 0.000 547.470 0.350 ;
    END
  END r0_rd_out[236]
  PIN r0_rd_out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 549.630 0.000 549.770 0.350 ;
    END
  END r0_rd_out[237]
  PIN r0_rd_out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 551.930 0.000 552.070 0.350 ;
    END
  END r0_rd_out[238]
  PIN r0_rd_out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 554.230 0.000 554.370 0.350 ;
    END
  END r0_rd_out[239]
  PIN r0_rd_out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 556.530 0.000 556.670 0.350 ;
    END
  END r0_rd_out[240]
  PIN r0_rd_out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 558.830 0.000 558.970 0.350 ;
    END
  END r0_rd_out[241]
  PIN r0_rd_out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 561.130 0.000 561.270 0.350 ;
    END
  END r0_rd_out[242]
  PIN r0_rd_out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 563.430 0.000 563.570 0.350 ;
    END
  END r0_rd_out[243]
  PIN r0_rd_out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 565.730 0.000 565.870 0.350 ;
    END
  END r0_rd_out[244]
  PIN r0_rd_out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 568.030 0.000 568.170 0.350 ;
    END
  END r0_rd_out[245]
  PIN r0_rd_out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 570.330 0.000 570.470 0.350 ;
    END
  END r0_rd_out[246]
  PIN r0_rd_out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 572.630 0.000 572.770 0.350 ;
    END
  END r0_rd_out[247]
  PIN r0_rd_out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 574.930 0.000 575.070 0.350 ;
    END
  END r0_rd_out[248]
  PIN r0_rd_out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 577.230 0.000 577.370 0.350 ;
    END
  END r0_rd_out[249]
  PIN r0_rd_out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 579.530 0.000 579.670 0.350 ;
    END
  END r0_rd_out[250]
  PIN r0_rd_out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 581.830 0.000 581.970 0.350 ;
    END
  END r0_rd_out[251]
  PIN r0_rd_out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 584.130 0.000 584.270 0.350 ;
    END
  END r0_rd_out[252]
  PIN r0_rd_out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 586.430 0.000 586.570 0.350 ;
    END
  END r0_rd_out[253]
  PIN r0_rd_out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 588.730 0.000 588.870 0.350 ;
    END
  END r0_rd_out[254]
  PIN r0_rd_out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 591.030 0.000 591.170 0.350 ;
    END
  END r0_rd_out[255]
  PIN r0_rd_out[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 593.330 0.000 593.470 0.350 ;
    END
  END r0_rd_out[256]
  PIN r0_rd_out[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 595.630 0.000 595.770 0.350 ;
    END
  END r0_rd_out[257]
  PIN r0_rd_out[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 597.930 0.000 598.070 0.350 ;
    END
  END r0_rd_out[258]
  PIN r0_rd_out[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 600.230 0.000 600.370 0.350 ;
    END
  END r0_rd_out[259]
  PIN r0_rd_out[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 602.530 0.000 602.670 0.350 ;
    END
  END r0_rd_out[260]
  PIN r0_rd_out[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 604.830 0.000 604.970 0.350 ;
    END
  END r0_rd_out[261]
  PIN r0_rd_out[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 607.130 0.000 607.270 0.350 ;
    END
  END r0_rd_out[262]
  PIN r0_rd_out[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 609.430 0.000 609.570 0.350 ;
    END
  END r0_rd_out[263]
  PIN r0_rd_out[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 611.730 0.000 611.870 0.350 ;
    END
  END r0_rd_out[264]
  PIN r0_rd_out[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 614.030 0.000 614.170 0.350 ;
    END
  END r0_rd_out[265]
  PIN r0_rd_out[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 616.330 0.000 616.470 0.350 ;
    END
  END r0_rd_out[266]
  PIN r0_rd_out[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 618.630 0.000 618.770 0.350 ;
    END
  END r0_rd_out[267]
  PIN r0_rd_out[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 620.930 0.000 621.070 0.350 ;
    END
  END r0_rd_out[268]
  PIN r0_rd_out[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 623.230 0.000 623.370 0.350 ;
    END
  END r0_rd_out[269]
  PIN r0_rd_out[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 625.530 0.000 625.670 0.350 ;
    END
  END r0_rd_out[270]
  PIN r0_rd_out[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 627.830 0.000 627.970 0.350 ;
    END
  END r0_rd_out[271]
  PIN r0_rd_out[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 630.130 0.000 630.270 0.350 ;
    END
  END r0_rd_out[272]
  PIN r0_rd_out[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 632.430 0.000 632.570 0.350 ;
    END
  END r0_rd_out[273]
  PIN r0_rd_out[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 634.730 0.000 634.870 0.350 ;
    END
  END r0_rd_out[274]
  PIN r0_rd_out[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 637.030 0.000 637.170 0.350 ;
    END
  END r0_rd_out[275]
  PIN r0_rd_out[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 639.330 0.000 639.470 0.350 ;
    END
  END r0_rd_out[276]
  PIN r0_rd_out[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 641.630 0.000 641.770 0.350 ;
    END
  END r0_rd_out[277]
  PIN r0_rd_out[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 643.930 0.000 644.070 0.350 ;
    END
  END r0_rd_out[278]
  PIN r0_rd_out[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 646.230 0.000 646.370 0.350 ;
    END
  END r0_rd_out[279]
  PIN r0_rd_out[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 648.530 0.000 648.670 0.350 ;
    END
  END r0_rd_out[280]
  PIN r0_rd_out[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 650.830 0.000 650.970 0.350 ;
    END
  END r0_rd_out[281]
  PIN r0_rd_out[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 653.130 0.000 653.270 0.350 ;
    END
  END r0_rd_out[282]
  PIN r0_rd_out[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 655.430 0.000 655.570 0.350 ;
    END
  END r0_rd_out[283]
  PIN r0_rd_out[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 657.730 0.000 657.870 0.350 ;
    END
  END r0_rd_out[284]
  PIN r0_rd_out[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 660.030 0.000 660.170 0.350 ;
    END
  END r0_rd_out[285]
  PIN r0_rd_out[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 662.330 0.000 662.470 0.350 ;
    END
  END r0_rd_out[286]
  PIN r0_rd_out[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 664.630 0.000 664.770 0.350 ;
    END
  END r0_rd_out[287]
  PIN r0_rd_out[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 666.930 0.000 667.070 0.350 ;
    END
  END r0_rd_out[288]
  PIN r0_rd_out[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 669.230 0.000 669.370 0.350 ;
    END
  END r0_rd_out[289]
  PIN r0_rd_out[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 671.530 0.000 671.670 0.350 ;
    END
  END r0_rd_out[290]
  PIN r0_rd_out[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 673.830 0.000 673.970 0.350 ;
    END
  END r0_rd_out[291]
  PIN r0_rd_out[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 676.130 0.000 676.270 0.350 ;
    END
  END r0_rd_out[292]
  PIN r0_rd_out[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 678.430 0.000 678.570 0.350 ;
    END
  END r0_rd_out[293]
  PIN r0_rd_out[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 680.730 0.000 680.870 0.350 ;
    END
  END r0_rd_out[294]
  PIN r0_rd_out[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 683.030 0.000 683.170 0.350 ;
    END
  END r0_rd_out[295]
  PIN r0_rd_out[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 685.330 0.000 685.470 0.350 ;
    END
  END r0_rd_out[296]
  PIN r0_rd_out[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 687.630 0.000 687.770 0.350 ;
    END
  END r0_rd_out[297]
  PIN r0_rd_out[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 689.930 0.000 690.070 0.350 ;
    END
  END r0_rd_out[298]
  PIN r0_rd_out[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 692.230 0.000 692.370 0.350 ;
    END
  END r0_rd_out[299]
  PIN r0_rd_out[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 694.530 0.000 694.670 0.350 ;
    END
  END r0_rd_out[300]
  PIN r0_rd_out[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 696.830 0.000 696.970 0.350 ;
    END
  END r0_rd_out[301]
  PIN r0_rd_out[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 699.130 0.000 699.270 0.350 ;
    END
  END r0_rd_out[302]
  PIN r0_rd_out[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 701.430 0.000 701.570 0.350 ;
    END
  END r0_rd_out[303]
  PIN r0_rd_out[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 703.730 0.000 703.870 0.350 ;
    END
  END r0_rd_out[304]
  PIN r0_rd_out[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 706.030 0.000 706.170 0.350 ;
    END
  END r0_rd_out[305]
  PIN r0_rd_out[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 708.330 0.000 708.470 0.350 ;
    END
  END r0_rd_out[306]
  PIN r0_rd_out[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 710.630 0.000 710.770 0.350 ;
    END
  END r0_rd_out[307]
  PIN r0_rd_out[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 712.930 0.000 713.070 0.350 ;
    END
  END r0_rd_out[308]
  PIN r0_rd_out[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 715.230 0.000 715.370 0.350 ;
    END
  END r0_rd_out[309]
  PIN r0_rd_out[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 717.530 0.000 717.670 0.350 ;
    END
  END r0_rd_out[310]
  PIN r0_rd_out[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 719.830 0.000 719.970 0.350 ;
    END
  END r0_rd_out[311]
  PIN r0_rd_out[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 722.130 0.000 722.270 0.350 ;
    END
  END r0_rd_out[312]
  PIN r0_rd_out[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 724.430 0.000 724.570 0.350 ;
    END
  END r0_rd_out[313]
  PIN r0_rd_out[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 726.730 0.000 726.870 0.350 ;
    END
  END r0_rd_out[314]
  PIN r0_rd_out[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 729.030 0.000 729.170 0.350 ;
    END
  END r0_rd_out[315]
  PIN r0_rd_out[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 731.330 0.000 731.470 0.350 ;
    END
  END r0_rd_out[316]
  PIN r0_rd_out[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 733.630 0.000 733.770 0.350 ;
    END
  END r0_rd_out[317]
  PIN r0_rd_out[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 735.930 0.000 736.070 0.350 ;
    END
  END r0_rd_out[318]
  PIN r0_rd_out[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 738.230 0.000 738.370 0.350 ;
    END
  END r0_rd_out[319]
  PIN r0_rd_out[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 740.530 0.000 740.670 0.350 ;
    END
  END r0_rd_out[320]
  PIN r0_rd_out[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 742.830 0.000 742.970 0.350 ;
    END
  END r0_rd_out[321]
  PIN r0_rd_out[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 745.130 0.000 745.270 0.350 ;
    END
  END r0_rd_out[322]
  PIN r0_rd_out[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 747.430 0.000 747.570 0.350 ;
    END
  END r0_rd_out[323]
  PIN r0_rd_out[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 749.730 0.000 749.870 0.350 ;
    END
  END r0_rd_out[324]
  PIN r0_rd_out[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 752.030 0.000 752.170 0.350 ;
    END
  END r0_rd_out[325]
  PIN r0_rd_out[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 754.330 0.000 754.470 0.350 ;
    END
  END r0_rd_out[326]
  PIN r0_rd_out[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 756.630 0.000 756.770 0.350 ;
    END
  END r0_rd_out[327]
  PIN r0_rd_out[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 758.930 0.000 759.070 0.350 ;
    END
  END r0_rd_out[328]
  PIN r0_rd_out[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 761.230 0.000 761.370 0.350 ;
    END
  END r0_rd_out[329]
  PIN r0_rd_out[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 763.530 0.000 763.670 0.350 ;
    END
  END r0_rd_out[330]
  PIN r0_rd_out[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 765.830 0.000 765.970 0.350 ;
    END
  END r0_rd_out[331]
  PIN r0_rd_out[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 768.130 0.000 768.270 0.350 ;
    END
  END r0_rd_out[332]
  PIN r0_rd_out[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 770.430 0.000 770.570 0.350 ;
    END
  END r0_rd_out[333]
  PIN r0_rd_out[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 772.730 0.000 772.870 0.350 ;
    END
  END r0_rd_out[334]
  PIN r0_rd_out[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 775.030 0.000 775.170 0.350 ;
    END
  END r0_rd_out[335]
  PIN r0_rd_out[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 777.330 0.000 777.470 0.350 ;
    END
  END r0_rd_out[336]
  PIN r0_rd_out[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 779.630 0.000 779.770 0.350 ;
    END
  END r0_rd_out[337]
  PIN r0_rd_out[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 781.930 0.000 782.070 0.350 ;
    END
  END r0_rd_out[338]
  PIN r0_rd_out[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 784.230 0.000 784.370 0.350 ;
    END
  END r0_rd_out[339]
  PIN r0_rd_out[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 786.530 0.000 786.670 0.350 ;
    END
  END r0_rd_out[340]
  PIN r0_rd_out[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 788.830 0.000 788.970 0.350 ;
    END
  END r0_rd_out[341]
  PIN r0_rd_out[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 791.130 0.000 791.270 0.350 ;
    END
  END r0_rd_out[342]
  PIN r0_rd_out[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 793.430 0.000 793.570 0.350 ;
    END
  END r0_rd_out[343]
  PIN r0_rd_out[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 795.730 0.000 795.870 0.350 ;
    END
  END r0_rd_out[344]
  PIN r0_rd_out[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 798.030 0.000 798.170 0.350 ;
    END
  END r0_rd_out[345]
  PIN r0_rd_out[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 800.330 0.000 800.470 0.350 ;
    END
  END r0_rd_out[346]
  PIN r0_rd_out[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 802.630 0.000 802.770 0.350 ;
    END
  END r0_rd_out[347]
  PIN r0_rd_out[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 804.930 0.000 805.070 0.350 ;
    END
  END r0_rd_out[348]
  PIN r0_rd_out[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 807.230 0.000 807.370 0.350 ;
    END
  END r0_rd_out[349]
  PIN r0_rd_out[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 809.530 0.000 809.670 0.350 ;
    END
  END r0_rd_out[350]
  PIN r0_rd_out[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 811.830 0.000 811.970 0.350 ;
    END
  END r0_rd_out[351]
  PIN r0_rd_out[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 814.130 0.000 814.270 0.350 ;
    END
  END r0_rd_out[352]
  PIN r0_rd_out[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 816.430 0.000 816.570 0.350 ;
    END
  END r0_rd_out[353]
  PIN r0_rd_out[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 818.730 0.000 818.870 0.350 ;
    END
  END r0_rd_out[354]
  PIN r0_rd_out[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 821.030 0.000 821.170 0.350 ;
    END
  END r0_rd_out[355]
  PIN r0_rd_out[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 823.330 0.000 823.470 0.350 ;
    END
  END r0_rd_out[356]
  PIN r0_rd_out[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 825.630 0.000 825.770 0.350 ;
    END
  END r0_rd_out[357]
  PIN r0_rd_out[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 827.930 0.000 828.070 0.350 ;
    END
  END r0_rd_out[358]
  PIN r0_rd_out[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 830.230 0.000 830.370 0.350 ;
    END
  END r0_rd_out[359]
  PIN r0_rd_out[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 832.530 0.000 832.670 0.350 ;
    END
  END r0_rd_out[360]
  PIN r0_rd_out[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 834.830 0.000 834.970 0.350 ;
    END
  END r0_rd_out[361]
  PIN r0_rd_out[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 837.130 0.000 837.270 0.350 ;
    END
  END r0_rd_out[362]
  PIN r0_rd_out[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 839.430 0.000 839.570 0.350 ;
    END
  END r0_rd_out[363]
  PIN r0_rd_out[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 841.730 0.000 841.870 0.350 ;
    END
  END r0_rd_out[364]
  PIN r0_rd_out[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 844.030 0.000 844.170 0.350 ;
    END
  END r0_rd_out[365]
  PIN r0_rd_out[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 846.330 0.000 846.470 0.350 ;
    END
  END r0_rd_out[366]
  PIN r0_rd_out[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 848.630 0.000 848.770 0.350 ;
    END
  END r0_rd_out[367]
  PIN r0_rd_out[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 850.930 0.000 851.070 0.350 ;
    END
  END r0_rd_out[368]
  PIN r0_rd_out[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 853.230 0.000 853.370 0.350 ;
    END
  END r0_rd_out[369]
  PIN r0_rd_out[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 855.530 0.000 855.670 0.350 ;
    END
  END r0_rd_out[370]
  PIN r0_rd_out[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 857.830 0.000 857.970 0.350 ;
    END
  END r0_rd_out[371]
  PIN r0_rd_out[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 860.130 0.000 860.270 0.350 ;
    END
  END r0_rd_out[372]
  PIN r0_rd_out[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 862.430 0.000 862.570 0.350 ;
    END
  END r0_rd_out[373]
  PIN r0_rd_out[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 864.730 0.000 864.870 0.350 ;
    END
  END r0_rd_out[374]
  PIN r0_rd_out[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 867.030 0.000 867.170 0.350 ;
    END
  END r0_rd_out[375]
  PIN r0_rd_out[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 869.330 0.000 869.470 0.350 ;
    END
  END r0_rd_out[376]
  PIN r0_rd_out[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 871.630 0.000 871.770 0.350 ;
    END
  END r0_rd_out[377]
  PIN r0_rd_out[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 873.930 0.000 874.070 0.350 ;
    END
  END r0_rd_out[378]
  PIN r0_rd_out[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 876.230 0.000 876.370 0.350 ;
    END
  END r0_rd_out[379]
  PIN r0_rd_out[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 878.530 0.000 878.670 0.350 ;
    END
  END r0_rd_out[380]
  PIN r0_rd_out[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 880.830 0.000 880.970 0.350 ;
    END
  END r0_rd_out[381]
  PIN r0_rd_out[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 883.130 0.000 883.270 0.350 ;
    END
  END r0_rd_out[382]
  PIN r0_rd_out[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 885.430 0.000 885.570 0.350 ;
    END
  END r0_rd_out[383]
  PIN r0_rd_out[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 887.730 0.000 887.870 0.350 ;
    END
  END r0_rd_out[384]
  PIN r0_rd_out[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 890.030 0.000 890.170 0.350 ;
    END
  END r0_rd_out[385]
  PIN r0_rd_out[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 892.330 0.000 892.470 0.350 ;
    END
  END r0_rd_out[386]
  PIN r0_rd_out[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 894.630 0.000 894.770 0.350 ;
    END
  END r0_rd_out[387]
  PIN r0_rd_out[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 896.930 0.000 897.070 0.350 ;
    END
  END r0_rd_out[388]
  PIN r0_rd_out[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 899.230 0.000 899.370 0.350 ;
    END
  END r0_rd_out[389]
  PIN r0_rd_out[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 901.530 0.000 901.670 0.350 ;
    END
  END r0_rd_out[390]
  PIN r0_rd_out[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 903.830 0.000 903.970 0.350 ;
    END
  END r0_rd_out[391]
  PIN r0_rd_out[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 906.130 0.000 906.270 0.350 ;
    END
  END r0_rd_out[392]
  PIN r0_rd_out[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 908.430 0.000 908.570 0.350 ;
    END
  END r0_rd_out[393]
  PIN r0_rd_out[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 910.730 0.000 910.870 0.350 ;
    END
  END r0_rd_out[394]
  PIN r0_rd_out[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 913.030 0.000 913.170 0.350 ;
    END
  END r0_rd_out[395]
  PIN r0_rd_out[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 915.330 0.000 915.470 0.350 ;
    END
  END r0_rd_out[396]
  PIN r0_rd_out[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 917.630 0.000 917.770 0.350 ;
    END
  END r0_rd_out[397]
  PIN r0_rd_out[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 919.930 0.000 920.070 0.350 ;
    END
  END r0_rd_out[398]
  PIN r0_rd_out[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 922.230 0.000 922.370 0.350 ;
    END
  END r0_rd_out[399]
  PIN r0_rd_out[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 924.530 0.000 924.670 0.350 ;
    END
  END r0_rd_out[400]
  PIN r0_rd_out[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 926.830 0.000 926.970 0.350 ;
    END
  END r0_rd_out[401]
  PIN r0_rd_out[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 929.130 0.000 929.270 0.350 ;
    END
  END r0_rd_out[402]
  PIN r0_rd_out[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 931.430 0.000 931.570 0.350 ;
    END
  END r0_rd_out[403]
  PIN r0_rd_out[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 933.730 0.000 933.870 0.350 ;
    END
  END r0_rd_out[404]
  PIN r0_rd_out[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 936.030 0.000 936.170 0.350 ;
    END
  END r0_rd_out[405]
  PIN r0_rd_out[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 938.330 0.000 938.470 0.350 ;
    END
  END r0_rd_out[406]
  PIN r0_rd_out[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 940.630 0.000 940.770 0.350 ;
    END
  END r0_rd_out[407]
  PIN r0_rd_out[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 942.930 0.000 943.070 0.350 ;
    END
  END r0_rd_out[408]
  PIN r0_rd_out[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 945.230 0.000 945.370 0.350 ;
    END
  END r0_rd_out[409]
  PIN r0_rd_out[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 947.530 0.000 947.670 0.350 ;
    END
  END r0_rd_out[410]
  PIN r0_rd_out[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 949.830 0.000 949.970 0.350 ;
    END
  END r0_rd_out[411]
  PIN r0_rd_out[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 952.130 0.000 952.270 0.350 ;
    END
  END r0_rd_out[412]
  PIN r0_rd_out[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 954.430 0.000 954.570 0.350 ;
    END
  END r0_rd_out[413]
  PIN r0_rd_out[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 956.730 0.000 956.870 0.350 ;
    END
  END r0_rd_out[414]
  PIN r0_rd_out[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 959.030 0.000 959.170 0.350 ;
    END
  END r0_rd_out[415]
  PIN r0_rd_out[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 961.330 0.000 961.470 0.350 ;
    END
  END r0_rd_out[416]
  PIN r0_rd_out[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 963.630 0.000 963.770 0.350 ;
    END
  END r0_rd_out[417]
  PIN r0_rd_out[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 965.930 0.000 966.070 0.350 ;
    END
  END r0_rd_out[418]
  PIN r0_rd_out[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 968.230 0.000 968.370 0.350 ;
    END
  END r0_rd_out[419]
  PIN r0_rd_out[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 970.530 0.000 970.670 0.350 ;
    END
  END r0_rd_out[420]
  PIN r0_rd_out[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 972.830 0.000 972.970 0.350 ;
    END
  END r0_rd_out[421]
  PIN r0_rd_out[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 975.130 0.000 975.270 0.350 ;
    END
  END r0_rd_out[422]
  PIN r0_rd_out[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 977.430 0.000 977.570 0.350 ;
    END
  END r0_rd_out[423]
  PIN r0_rd_out[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 979.730 0.000 979.870 0.350 ;
    END
  END r0_rd_out[424]
  PIN r0_rd_out[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 982.030 0.000 982.170 0.350 ;
    END
  END r0_rd_out[425]
  PIN r0_rd_out[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 984.330 0.000 984.470 0.350 ;
    END
  END r0_rd_out[426]
  PIN r0_rd_out[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 986.630 0.000 986.770 0.350 ;
    END
  END r0_rd_out[427]
  PIN r0_rd_out[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 988.930 0.000 989.070 0.350 ;
    END
  END r0_rd_out[428]
  PIN r0_rd_out[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 991.230 0.000 991.370 0.350 ;
    END
  END r0_rd_out[429]
  PIN r0_rd_out[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 993.530 0.000 993.670 0.350 ;
    END
  END r0_rd_out[430]
  PIN r0_rd_out[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 995.830 0.000 995.970 0.350 ;
    END
  END r0_rd_out[431]
  PIN r0_rd_out[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 998.130 0.000 998.270 0.350 ;
    END
  END r0_rd_out[432]
  PIN r0_rd_out[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1000.430 0.000 1000.570 0.350 ;
    END
  END r0_rd_out[433]
  PIN r0_rd_out[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1002.730 0.000 1002.870 0.350 ;
    END
  END r0_rd_out[434]
  PIN r0_rd_out[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1005.030 0.000 1005.170 0.350 ;
    END
  END r0_rd_out[435]
  PIN r0_rd_out[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1007.330 0.000 1007.470 0.350 ;
    END
  END r0_rd_out[436]
  PIN r0_rd_out[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1009.630 0.000 1009.770 0.350 ;
    END
  END r0_rd_out[437]
  PIN r0_rd_out[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1011.930 0.000 1012.070 0.350 ;
    END
  END r0_rd_out[438]
  PIN r0_rd_out[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1014.230 0.000 1014.370 0.350 ;
    END
  END r0_rd_out[439]
  PIN r0_rd_out[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1016.530 0.000 1016.670 0.350 ;
    END
  END r0_rd_out[440]
  PIN r0_rd_out[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1018.830 0.000 1018.970 0.350 ;
    END
  END r0_rd_out[441]
  PIN r0_rd_out[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1021.130 0.000 1021.270 0.350 ;
    END
  END r0_rd_out[442]
  PIN r0_rd_out[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1023.430 0.000 1023.570 0.350 ;
    END
  END r0_rd_out[443]
  PIN r0_rd_out[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1025.730 0.000 1025.870 0.350 ;
    END
  END r0_rd_out[444]
  PIN r0_rd_out[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1028.030 0.000 1028.170 0.350 ;
    END
  END r0_rd_out[445]
  PIN r0_rd_out[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1030.330 0.000 1030.470 0.350 ;
    END
  END r0_rd_out[446]
  PIN r0_rd_out[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1032.630 0.000 1032.770 0.350 ;
    END
  END r0_rd_out[447]
  PIN r0_rd_out[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1034.930 0.000 1035.070 0.350 ;
    END
  END r0_rd_out[448]
  PIN r0_rd_out[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1037.230 0.000 1037.370 0.350 ;
    END
  END r0_rd_out[449]
  PIN r0_rd_out[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1039.530 0.000 1039.670 0.350 ;
    END
  END r0_rd_out[450]
  PIN r0_rd_out[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1041.830 0.000 1041.970 0.350 ;
    END
  END r0_rd_out[451]
  PIN r0_rd_out[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1044.130 0.000 1044.270 0.350 ;
    END
  END r0_rd_out[452]
  PIN r0_rd_out[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1046.430 0.000 1046.570 0.350 ;
    END
  END r0_rd_out[453]
  PIN r0_rd_out[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1048.730 0.000 1048.870 0.350 ;
    END
  END r0_rd_out[454]
  PIN r0_rd_out[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1051.030 0.000 1051.170 0.350 ;
    END
  END r0_rd_out[455]
  PIN r0_rd_out[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1053.330 0.000 1053.470 0.350 ;
    END
  END r0_rd_out[456]
  PIN r0_rd_out[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1055.630 0.000 1055.770 0.350 ;
    END
  END r0_rd_out[457]
  PIN r0_rd_out[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1057.930 0.000 1058.070 0.350 ;
    END
  END r0_rd_out[458]
  PIN r0_rd_out[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1060.230 0.000 1060.370 0.350 ;
    END
  END r0_rd_out[459]
  PIN r0_rd_out[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1062.530 0.000 1062.670 0.350 ;
    END
  END r0_rd_out[460]
  PIN r0_rd_out[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1064.830 0.000 1064.970 0.350 ;
    END
  END r0_rd_out[461]
  PIN r0_rd_out[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1067.130 0.000 1067.270 0.350 ;
    END
  END r0_rd_out[462]
  PIN r0_rd_out[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1069.430 0.000 1069.570 0.350 ;
    END
  END r0_rd_out[463]
  PIN r0_rd_out[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1071.730 0.000 1071.870 0.350 ;
    END
  END r0_rd_out[464]
  PIN r0_rd_out[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1074.030 0.000 1074.170 0.350 ;
    END
  END r0_rd_out[465]
  PIN r0_rd_out[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1076.330 0.000 1076.470 0.350 ;
    END
  END r0_rd_out[466]
  PIN r0_rd_out[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1078.630 0.000 1078.770 0.350 ;
    END
  END r0_rd_out[467]
  PIN r0_rd_out[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1080.930 0.000 1081.070 0.350 ;
    END
  END r0_rd_out[468]
  PIN r0_rd_out[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1083.230 0.000 1083.370 0.350 ;
    END
  END r0_rd_out[469]
  PIN r0_rd_out[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1085.530 0.000 1085.670 0.350 ;
    END
  END r0_rd_out[470]
  PIN r0_rd_out[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1087.830 0.000 1087.970 0.350 ;
    END
  END r0_rd_out[471]
  PIN r0_rd_out[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1090.130 0.000 1090.270 0.350 ;
    END
  END r0_rd_out[472]
  PIN r0_rd_out[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1092.430 0.000 1092.570 0.350 ;
    END
  END r0_rd_out[473]
  PIN r0_rd_out[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1094.730 0.000 1094.870 0.350 ;
    END
  END r0_rd_out[474]
  PIN r0_rd_out[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1097.030 0.000 1097.170 0.350 ;
    END
  END r0_rd_out[475]
  PIN r0_rd_out[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1099.330 0.000 1099.470 0.350 ;
    END
  END r0_rd_out[476]
  PIN r0_rd_out[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1101.630 0.000 1101.770 0.350 ;
    END
  END r0_rd_out[477]
  PIN r0_rd_out[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1103.930 0.000 1104.070 0.350 ;
    END
  END r0_rd_out[478]
  PIN r0_rd_out[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1106.230 0.000 1106.370 0.350 ;
    END
  END r0_rd_out[479]
  PIN r0_rd_out[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1108.530 0.000 1108.670 0.350 ;
    END
  END r0_rd_out[480]
  PIN r0_rd_out[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1110.830 0.000 1110.970 0.350 ;
    END
  END r0_rd_out[481]
  PIN r0_rd_out[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1113.130 0.000 1113.270 0.350 ;
    END
  END r0_rd_out[482]
  PIN r0_rd_out[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1115.430 0.000 1115.570 0.350 ;
    END
  END r0_rd_out[483]
  PIN r0_rd_out[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1117.730 0.000 1117.870 0.350 ;
    END
  END r0_rd_out[484]
  PIN r0_rd_out[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1120.030 0.000 1120.170 0.350 ;
    END
  END r0_rd_out[485]
  PIN r0_rd_out[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1122.330 0.000 1122.470 0.350 ;
    END
  END r0_rd_out[486]
  PIN r0_rd_out[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1124.630 0.000 1124.770 0.350 ;
    END
  END r0_rd_out[487]
  PIN r0_rd_out[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1126.930 0.000 1127.070 0.350 ;
    END
  END r0_rd_out[488]
  PIN r0_rd_out[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1129.230 0.000 1129.370 0.350 ;
    END
  END r0_rd_out[489]
  PIN r0_rd_out[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1131.530 0.000 1131.670 0.350 ;
    END
  END r0_rd_out[490]
  PIN r0_rd_out[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1133.830 0.000 1133.970 0.350 ;
    END
  END r0_rd_out[491]
  PIN r0_rd_out[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1136.130 0.000 1136.270 0.350 ;
    END
  END r0_rd_out[492]
  PIN r0_rd_out[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1138.430 0.000 1138.570 0.350 ;
    END
  END r0_rd_out[493]
  PIN r0_rd_out[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1140.730 0.000 1140.870 0.350 ;
    END
  END r0_rd_out[494]
  PIN r0_rd_out[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1143.030 0.000 1143.170 0.350 ;
    END
  END r0_rd_out[495]
  PIN r0_rd_out[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1145.330 0.000 1145.470 0.350 ;
    END
  END r0_rd_out[496]
  PIN r0_rd_out[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1147.630 0.000 1147.770 0.350 ;
    END
  END r0_rd_out[497]
  PIN r0_rd_out[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1149.930 0.000 1150.070 0.350 ;
    END
  END r0_rd_out[498]
  PIN r0_rd_out[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1152.230 0.000 1152.370 0.350 ;
    END
  END r0_rd_out[499]
  PIN r0_rd_out[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1154.530 0.000 1154.670 0.350 ;
    END
  END r0_rd_out[500]
  PIN r0_rd_out[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1156.830 0.000 1156.970 0.350 ;
    END
  END r0_rd_out[501]
  PIN r0_rd_out[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1159.130 0.000 1159.270 0.350 ;
    END
  END r0_rd_out[502]
  PIN r0_rd_out[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1161.430 0.000 1161.570 0.350 ;
    END
  END r0_rd_out[503]
  PIN r0_rd_out[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1163.730 0.000 1163.870 0.350 ;
    END
  END r0_rd_out[504]
  PIN r0_rd_out[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1166.030 0.000 1166.170 0.350 ;
    END
  END r0_rd_out[505]
  PIN r0_rd_out[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1168.330 0.000 1168.470 0.350 ;
    END
  END r0_rd_out[506]
  PIN r0_rd_out[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1170.630 0.000 1170.770 0.350 ;
    END
  END r0_rd_out[507]
  PIN r0_rd_out[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1172.930 0.000 1173.070 0.350 ;
    END
  END r0_rd_out[508]
  PIN r0_rd_out[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1175.230 0.000 1175.370 0.350 ;
    END
  END r0_rd_out[509]
  PIN r0_rd_out[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1177.530 0.000 1177.670 0.350 ;
    END
  END r0_rd_out[510]
  PIN r0_rd_out[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 1179.830 0.000 1179.970 0.350 ;
    END
  END r0_rd_out[511]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 1301.920 6.650 1302.720 6.950 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 1301.920 9.370 1302.720 9.670 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 1301.920 12.090 1302.720 12.390 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 1301.920 14.810 1302.720 15.110 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 1301.920 17.530 1302.720 17.830 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 1301.920 20.250 1302.720 20.550 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 1301.920 22.970 1302.720 23.270 ;
    END
  END w0_addr_in[6]
  PIN w0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 1301.920 25.690 1302.720 25.990 ;
    END
  END w0_addr_in[7]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 4.530 1569.090 4.670 1569.440 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 6.830 1569.090 6.970 1569.440 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 9.130 1569.090 9.270 1569.440 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 11.430 1569.090 11.570 1569.440 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 13.730 1569.090 13.870 1569.440 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 16.030 1569.090 16.170 1569.440 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 18.330 1569.090 18.470 1569.440 ;
    END
  END r0_addr_in[6]
  PIN r0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 20.630 1569.090 20.770 1569.440 ;
    END
  END r0_addr_in[7]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 1301.920 103.210 1302.720 103.510 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 1301.920 180.730 1302.720 181.030 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 1301.920 258.250 1302.720 258.550 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 76.290 1569.090 76.430 1569.440 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
      RECT 131.950 1569.090 132.090 1569.440 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 3.240 6.800 5.960 1562.640 ;
      RECT 14.120 6.800 16.840 1562.640 ;
      RECT 25.000 6.800 27.720 1562.640 ;
      RECT 35.880 6.800 38.600 1562.640 ;
      RECT 46.760 6.800 49.480 1562.640 ;
      RECT 57.640 6.800 60.360 1562.640 ;
      RECT 68.520 6.800 71.240 1562.640 ;
      RECT 79.400 6.800 82.120 1562.640 ;
      RECT 90.280 6.800 93.000 1562.640 ;
      RECT 101.160 6.800 103.880 1562.640 ;
      RECT 112.040 6.800 114.760 1562.640 ;
      RECT 122.920 6.800 125.640 1562.640 ;
      RECT 133.800 6.800 136.520 1562.640 ;
      RECT 144.680 6.800 147.400 1562.640 ;
      RECT 155.560 6.800 158.280 1562.640 ;
      RECT 166.440 6.800 169.160 1562.640 ;
      RECT 177.320 6.800 180.040 1562.640 ;
      RECT 188.200 6.800 190.920 1562.640 ;
      RECT 199.080 6.800 201.800 1562.640 ;
      RECT 209.960 6.800 212.680 1562.640 ;
      RECT 220.840 6.800 223.560 1562.640 ;
      RECT 231.720 6.800 234.440 1562.640 ;
      RECT 242.600 6.800 245.320 1562.640 ;
      RECT 253.480 6.800 256.200 1562.640 ;
      RECT 264.360 6.800 267.080 1562.640 ;
      RECT 275.240 6.800 277.960 1562.640 ;
      RECT 286.120 6.800 288.840 1562.640 ;
      RECT 297.000 6.800 299.720 1562.640 ;
      RECT 307.880 6.800 310.600 1562.640 ;
      RECT 318.760 6.800 321.480 1562.640 ;
      RECT 329.640 6.800 332.360 1562.640 ;
      RECT 340.520 6.800 343.240 1562.640 ;
      RECT 351.400 6.800 354.120 1562.640 ;
      RECT 362.280 6.800 365.000 1562.640 ;
      RECT 373.160 6.800 375.880 1562.640 ;
      RECT 384.040 6.800 386.760 1562.640 ;
      RECT 394.920 6.800 397.640 1562.640 ;
      RECT 405.800 6.800 408.520 1562.640 ;
      RECT 416.680 6.800 419.400 1562.640 ;
      RECT 427.560 6.800 430.280 1562.640 ;
      RECT 438.440 6.800 441.160 1562.640 ;
      RECT 449.320 6.800 452.040 1562.640 ;
      RECT 460.200 6.800 462.920 1562.640 ;
      RECT 471.080 6.800 473.800 1562.640 ;
      RECT 481.960 6.800 484.680 1562.640 ;
      RECT 492.840 6.800 495.560 1562.640 ;
      RECT 503.720 6.800 506.440 1562.640 ;
      RECT 514.600 6.800 517.320 1562.640 ;
      RECT 525.480 6.800 528.200 1562.640 ;
      RECT 536.360 6.800 539.080 1562.640 ;
      RECT 547.240 6.800 549.960 1562.640 ;
      RECT 558.120 6.800 560.840 1562.640 ;
      RECT 569.000 6.800 571.720 1562.640 ;
      RECT 579.880 6.800 582.600 1562.640 ;
      RECT 590.760 6.800 593.480 1562.640 ;
      RECT 601.640 6.800 604.360 1562.640 ;
      RECT 612.520 6.800 615.240 1562.640 ;
      RECT 623.400 6.800 626.120 1562.640 ;
      RECT 634.280 6.800 637.000 1562.640 ;
      RECT 645.160 6.800 647.880 1562.640 ;
      RECT 656.040 6.800 658.760 1562.640 ;
      RECT 666.920 6.800 669.640 1562.640 ;
      RECT 677.800 6.800 680.520 1562.640 ;
      RECT 688.680 6.800 691.400 1562.640 ;
      RECT 699.560 6.800 702.280 1562.640 ;
      RECT 710.440 6.800 713.160 1562.640 ;
      RECT 721.320 6.800 724.040 1562.640 ;
      RECT 732.200 6.800 734.920 1562.640 ;
      RECT 743.080 6.800 745.800 1562.640 ;
      RECT 753.960 6.800 756.680 1562.640 ;
      RECT 764.840 6.800 767.560 1562.640 ;
      RECT 775.720 6.800 778.440 1562.640 ;
      RECT 786.600 6.800 789.320 1562.640 ;
      RECT 797.480 6.800 800.200 1562.640 ;
      RECT 808.360 6.800 811.080 1562.640 ;
      RECT 819.240 6.800 821.960 1562.640 ;
      RECT 830.120 6.800 832.840 1562.640 ;
      RECT 841.000 6.800 843.720 1562.640 ;
      RECT 851.880 6.800 854.600 1562.640 ;
      RECT 862.760 6.800 865.480 1562.640 ;
      RECT 873.640 6.800 876.360 1562.640 ;
      RECT 884.520 6.800 887.240 1562.640 ;
      RECT 895.400 6.800 898.120 1562.640 ;
      RECT 906.280 6.800 909.000 1562.640 ;
      RECT 917.160 6.800 919.880 1562.640 ;
      RECT 928.040 6.800 930.760 1562.640 ;
      RECT 938.920 6.800 941.640 1562.640 ;
      RECT 949.800 6.800 952.520 1562.640 ;
      RECT 960.680 6.800 963.400 1562.640 ;
      RECT 971.560 6.800 974.280 1562.640 ;
      RECT 982.440 6.800 985.160 1562.640 ;
      RECT 993.320 6.800 996.040 1562.640 ;
      RECT 1004.200 6.800 1006.920 1562.640 ;
      RECT 1015.080 6.800 1017.800 1562.640 ;
      RECT 1025.960 6.800 1028.680 1562.640 ;
      RECT 1036.840 6.800 1039.560 1562.640 ;
      RECT 1047.720 6.800 1050.440 1562.640 ;
      RECT 1058.600 6.800 1061.320 1562.640 ;
      RECT 1069.480 6.800 1072.200 1562.640 ;
      RECT 1080.360 6.800 1083.080 1562.640 ;
      RECT 1091.240 6.800 1093.960 1562.640 ;
      RECT 1102.120 6.800 1104.840 1562.640 ;
      RECT 1113.000 6.800 1115.720 1562.640 ;
      RECT 1123.880 6.800 1126.600 1562.640 ;
      RECT 1134.760 6.800 1137.480 1562.640 ;
      RECT 1145.640 6.800 1148.360 1562.640 ;
      RECT 1156.520 6.800 1159.240 1562.640 ;
      RECT 1167.400 6.800 1170.120 1562.640 ;
      RECT 1178.280 6.800 1181.000 1562.640 ;
      RECT 1189.160 6.800 1191.880 1562.640 ;
      RECT 1200.040 6.800 1202.760 1562.640 ;
      RECT 1210.920 6.800 1213.640 1562.640 ;
      RECT 1221.800 6.800 1224.520 1562.640 ;
      RECT 1232.680 6.800 1235.400 1562.640 ;
      RECT 1243.560 6.800 1246.280 1562.640 ;
      RECT 1254.440 6.800 1257.160 1562.640 ;
      RECT 1265.320 6.800 1268.040 1562.640 ;
      RECT 1276.200 6.800 1278.920 1562.640 ;
      RECT 1287.080 6.800 1289.800 1562.640 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 8.680 6.800 11.400 1562.640 ;
      RECT 19.560 6.800 22.280 1562.640 ;
      RECT 30.440 6.800 33.160 1562.640 ;
      RECT 41.320 6.800 44.040 1562.640 ;
      RECT 52.200 6.800 54.920 1562.640 ;
      RECT 63.080 6.800 65.800 1562.640 ;
      RECT 73.960 6.800 76.680 1562.640 ;
      RECT 84.840 6.800 87.560 1562.640 ;
      RECT 95.720 6.800 98.440 1562.640 ;
      RECT 106.600 6.800 109.320 1562.640 ;
      RECT 117.480 6.800 120.200 1562.640 ;
      RECT 128.360 6.800 131.080 1562.640 ;
      RECT 139.240 6.800 141.960 1562.640 ;
      RECT 150.120 6.800 152.840 1562.640 ;
      RECT 161.000 6.800 163.720 1562.640 ;
      RECT 171.880 6.800 174.600 1562.640 ;
      RECT 182.760 6.800 185.480 1562.640 ;
      RECT 193.640 6.800 196.360 1562.640 ;
      RECT 204.520 6.800 207.240 1562.640 ;
      RECT 215.400 6.800 218.120 1562.640 ;
      RECT 226.280 6.800 229.000 1562.640 ;
      RECT 237.160 6.800 239.880 1562.640 ;
      RECT 248.040 6.800 250.760 1562.640 ;
      RECT 258.920 6.800 261.640 1562.640 ;
      RECT 269.800 6.800 272.520 1562.640 ;
      RECT 280.680 6.800 283.400 1562.640 ;
      RECT 291.560 6.800 294.280 1562.640 ;
      RECT 302.440 6.800 305.160 1562.640 ;
      RECT 313.320 6.800 316.040 1562.640 ;
      RECT 324.200 6.800 326.920 1562.640 ;
      RECT 335.080 6.800 337.800 1562.640 ;
      RECT 345.960 6.800 348.680 1562.640 ;
      RECT 356.840 6.800 359.560 1562.640 ;
      RECT 367.720 6.800 370.440 1562.640 ;
      RECT 378.600 6.800 381.320 1562.640 ;
      RECT 389.480 6.800 392.200 1562.640 ;
      RECT 400.360 6.800 403.080 1562.640 ;
      RECT 411.240 6.800 413.960 1562.640 ;
      RECT 422.120 6.800 424.840 1562.640 ;
      RECT 433.000 6.800 435.720 1562.640 ;
      RECT 443.880 6.800 446.600 1562.640 ;
      RECT 454.760 6.800 457.480 1562.640 ;
      RECT 465.640 6.800 468.360 1562.640 ;
      RECT 476.520 6.800 479.240 1562.640 ;
      RECT 487.400 6.800 490.120 1562.640 ;
      RECT 498.280 6.800 501.000 1562.640 ;
      RECT 509.160 6.800 511.880 1562.640 ;
      RECT 520.040 6.800 522.760 1562.640 ;
      RECT 530.920 6.800 533.640 1562.640 ;
      RECT 541.800 6.800 544.520 1562.640 ;
      RECT 552.680 6.800 555.400 1562.640 ;
      RECT 563.560 6.800 566.280 1562.640 ;
      RECT 574.440 6.800 577.160 1562.640 ;
      RECT 585.320 6.800 588.040 1562.640 ;
      RECT 596.200 6.800 598.920 1562.640 ;
      RECT 607.080 6.800 609.800 1562.640 ;
      RECT 617.960 6.800 620.680 1562.640 ;
      RECT 628.840 6.800 631.560 1562.640 ;
      RECT 639.720 6.800 642.440 1562.640 ;
      RECT 650.600 6.800 653.320 1562.640 ;
      RECT 661.480 6.800 664.200 1562.640 ;
      RECT 672.360 6.800 675.080 1562.640 ;
      RECT 683.240 6.800 685.960 1562.640 ;
      RECT 694.120 6.800 696.840 1562.640 ;
      RECT 705.000 6.800 707.720 1562.640 ;
      RECT 715.880 6.800 718.600 1562.640 ;
      RECT 726.760 6.800 729.480 1562.640 ;
      RECT 737.640 6.800 740.360 1562.640 ;
      RECT 748.520 6.800 751.240 1562.640 ;
      RECT 759.400 6.800 762.120 1562.640 ;
      RECT 770.280 6.800 773.000 1562.640 ;
      RECT 781.160 6.800 783.880 1562.640 ;
      RECT 792.040 6.800 794.760 1562.640 ;
      RECT 802.920 6.800 805.640 1562.640 ;
      RECT 813.800 6.800 816.520 1562.640 ;
      RECT 824.680 6.800 827.400 1562.640 ;
      RECT 835.560 6.800 838.280 1562.640 ;
      RECT 846.440 6.800 849.160 1562.640 ;
      RECT 857.320 6.800 860.040 1562.640 ;
      RECT 868.200 6.800 870.920 1562.640 ;
      RECT 879.080 6.800 881.800 1562.640 ;
      RECT 889.960 6.800 892.680 1562.640 ;
      RECT 900.840 6.800 903.560 1562.640 ;
      RECT 911.720 6.800 914.440 1562.640 ;
      RECT 922.600 6.800 925.320 1562.640 ;
      RECT 933.480 6.800 936.200 1562.640 ;
      RECT 944.360 6.800 947.080 1562.640 ;
      RECT 955.240 6.800 957.960 1562.640 ;
      RECT 966.120 6.800 968.840 1562.640 ;
      RECT 977.000 6.800 979.720 1562.640 ;
      RECT 987.880 6.800 990.600 1562.640 ;
      RECT 998.760 6.800 1001.480 1562.640 ;
      RECT 1009.640 6.800 1012.360 1562.640 ;
      RECT 1020.520 6.800 1023.240 1562.640 ;
      RECT 1031.400 6.800 1034.120 1562.640 ;
      RECT 1042.280 6.800 1045.000 1562.640 ;
      RECT 1053.160 6.800 1055.880 1562.640 ;
      RECT 1064.040 6.800 1066.760 1562.640 ;
      RECT 1074.920 6.800 1077.640 1562.640 ;
      RECT 1085.800 6.800 1088.520 1562.640 ;
      RECT 1096.680 6.800 1099.400 1562.640 ;
      RECT 1107.560 6.800 1110.280 1562.640 ;
      RECT 1118.440 6.800 1121.160 1562.640 ;
      RECT 1129.320 6.800 1132.040 1562.640 ;
      RECT 1140.200 6.800 1142.920 1562.640 ;
      RECT 1151.080 6.800 1153.800 1562.640 ;
      RECT 1161.960 6.800 1164.680 1562.640 ;
      RECT 1172.840 6.800 1175.560 1562.640 ;
      RECT 1183.720 6.800 1186.440 1562.640 ;
      RECT 1194.600 6.800 1197.320 1562.640 ;
      RECT 1205.480 6.800 1208.200 1562.640 ;
      RECT 1216.360 6.800 1219.080 1562.640 ;
      RECT 1227.240 6.800 1229.960 1562.640 ;
      RECT 1238.120 6.800 1240.840 1562.640 ;
      RECT 1249.000 6.800 1251.720 1562.640 ;
      RECT 1259.880 6.800 1262.600 1562.640 ;
      RECT 1270.760 6.800 1273.480 1562.640 ;
      RECT 1281.640 6.800 1284.360 1562.640 ;
      RECT 1292.520 6.800 1295.240 1562.640 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 1302.720 1569.440 ;
    LAYER met2 ;
    RECT 0 0 1302.720 1569.440 ;
    LAYER met3 ;
    RECT 0.800 0 1302.720 1569.440 ;
    LAYER met4 ;
    RECT 0 0 1302.720 6.800 ;
    RECT 0 1562.640 1302.720 1569.440 ;
    RECT 0.000 6.800 3.240 1562.640 ;
    RECT 5.960 6.800 8.680 1562.640 ;
    RECT 11.400 6.800 14.120 1562.640 ;
    RECT 16.840 6.800 19.560 1562.640 ;
    RECT 22.280 6.800 25.000 1562.640 ;
    RECT 27.720 6.800 30.440 1562.640 ;
    RECT 33.160 6.800 35.880 1562.640 ;
    RECT 38.600 6.800 41.320 1562.640 ;
    RECT 44.040 6.800 46.760 1562.640 ;
    RECT 49.480 6.800 52.200 1562.640 ;
    RECT 54.920 6.800 57.640 1562.640 ;
    RECT 60.360 6.800 63.080 1562.640 ;
    RECT 65.800 6.800 68.520 1562.640 ;
    RECT 71.240 6.800 73.960 1562.640 ;
    RECT 76.680 6.800 79.400 1562.640 ;
    RECT 82.120 6.800 84.840 1562.640 ;
    RECT 87.560 6.800 90.280 1562.640 ;
    RECT 93.000 6.800 95.720 1562.640 ;
    RECT 98.440 6.800 101.160 1562.640 ;
    RECT 103.880 6.800 106.600 1562.640 ;
    RECT 109.320 6.800 112.040 1562.640 ;
    RECT 114.760 6.800 117.480 1562.640 ;
    RECT 120.200 6.800 122.920 1562.640 ;
    RECT 125.640 6.800 128.360 1562.640 ;
    RECT 131.080 6.800 133.800 1562.640 ;
    RECT 136.520 6.800 139.240 1562.640 ;
    RECT 141.960 6.800 144.680 1562.640 ;
    RECT 147.400 6.800 150.120 1562.640 ;
    RECT 152.840 6.800 155.560 1562.640 ;
    RECT 158.280 6.800 161.000 1562.640 ;
    RECT 163.720 6.800 166.440 1562.640 ;
    RECT 169.160 6.800 171.880 1562.640 ;
    RECT 174.600 6.800 177.320 1562.640 ;
    RECT 180.040 6.800 182.760 1562.640 ;
    RECT 185.480 6.800 188.200 1562.640 ;
    RECT 190.920 6.800 193.640 1562.640 ;
    RECT 196.360 6.800 199.080 1562.640 ;
    RECT 201.800 6.800 204.520 1562.640 ;
    RECT 207.240 6.800 209.960 1562.640 ;
    RECT 212.680 6.800 215.400 1562.640 ;
    RECT 218.120 6.800 220.840 1562.640 ;
    RECT 223.560 6.800 226.280 1562.640 ;
    RECT 229.000 6.800 231.720 1562.640 ;
    RECT 234.440 6.800 237.160 1562.640 ;
    RECT 239.880 6.800 242.600 1562.640 ;
    RECT 245.320 6.800 248.040 1562.640 ;
    RECT 250.760 6.800 253.480 1562.640 ;
    RECT 256.200 6.800 258.920 1562.640 ;
    RECT 261.640 6.800 264.360 1562.640 ;
    RECT 267.080 6.800 269.800 1562.640 ;
    RECT 272.520 6.800 275.240 1562.640 ;
    RECT 277.960 6.800 280.680 1562.640 ;
    RECT 283.400 6.800 286.120 1562.640 ;
    RECT 288.840 6.800 291.560 1562.640 ;
    RECT 294.280 6.800 297.000 1562.640 ;
    RECT 299.720 6.800 302.440 1562.640 ;
    RECT 305.160 6.800 307.880 1562.640 ;
    RECT 310.600 6.800 313.320 1562.640 ;
    RECT 316.040 6.800 318.760 1562.640 ;
    RECT 321.480 6.800 324.200 1562.640 ;
    RECT 326.920 6.800 329.640 1562.640 ;
    RECT 332.360 6.800 335.080 1562.640 ;
    RECT 337.800 6.800 340.520 1562.640 ;
    RECT 343.240 6.800 345.960 1562.640 ;
    RECT 348.680 6.800 351.400 1562.640 ;
    RECT 354.120 6.800 356.840 1562.640 ;
    RECT 359.560 6.800 362.280 1562.640 ;
    RECT 365.000 6.800 367.720 1562.640 ;
    RECT 370.440 6.800 373.160 1562.640 ;
    RECT 375.880 6.800 378.600 1562.640 ;
    RECT 381.320 6.800 384.040 1562.640 ;
    RECT 386.760 6.800 389.480 1562.640 ;
    RECT 392.200 6.800 394.920 1562.640 ;
    RECT 397.640 6.800 400.360 1562.640 ;
    RECT 403.080 6.800 405.800 1562.640 ;
    RECT 408.520 6.800 411.240 1562.640 ;
    RECT 413.960 6.800 416.680 1562.640 ;
    RECT 419.400 6.800 422.120 1562.640 ;
    RECT 424.840 6.800 427.560 1562.640 ;
    RECT 430.280 6.800 433.000 1562.640 ;
    RECT 435.720 6.800 438.440 1562.640 ;
    RECT 441.160 6.800 443.880 1562.640 ;
    RECT 446.600 6.800 449.320 1562.640 ;
    RECT 452.040 6.800 454.760 1562.640 ;
    RECT 457.480 6.800 460.200 1562.640 ;
    RECT 462.920 6.800 465.640 1562.640 ;
    RECT 468.360 6.800 471.080 1562.640 ;
    RECT 473.800 6.800 476.520 1562.640 ;
    RECT 479.240 6.800 481.960 1562.640 ;
    RECT 484.680 6.800 487.400 1562.640 ;
    RECT 490.120 6.800 492.840 1562.640 ;
    RECT 495.560 6.800 498.280 1562.640 ;
    RECT 501.000 6.800 503.720 1562.640 ;
    RECT 506.440 6.800 509.160 1562.640 ;
    RECT 511.880 6.800 514.600 1562.640 ;
    RECT 517.320 6.800 520.040 1562.640 ;
    RECT 522.760 6.800 525.480 1562.640 ;
    RECT 528.200 6.800 530.920 1562.640 ;
    RECT 533.640 6.800 536.360 1562.640 ;
    RECT 539.080 6.800 541.800 1562.640 ;
    RECT 544.520 6.800 547.240 1562.640 ;
    RECT 549.960 6.800 552.680 1562.640 ;
    RECT 555.400 6.800 558.120 1562.640 ;
    RECT 560.840 6.800 563.560 1562.640 ;
    RECT 566.280 6.800 569.000 1562.640 ;
    RECT 571.720 6.800 574.440 1562.640 ;
    RECT 577.160 6.800 579.880 1562.640 ;
    RECT 582.600 6.800 585.320 1562.640 ;
    RECT 588.040 6.800 590.760 1562.640 ;
    RECT 593.480 6.800 596.200 1562.640 ;
    RECT 598.920 6.800 601.640 1562.640 ;
    RECT 604.360 6.800 607.080 1562.640 ;
    RECT 609.800 6.800 612.520 1562.640 ;
    RECT 615.240 6.800 617.960 1562.640 ;
    RECT 620.680 6.800 623.400 1562.640 ;
    RECT 626.120 6.800 628.840 1562.640 ;
    RECT 631.560 6.800 634.280 1562.640 ;
    RECT 637.000 6.800 639.720 1562.640 ;
    RECT 642.440 6.800 645.160 1562.640 ;
    RECT 647.880 6.800 650.600 1562.640 ;
    RECT 653.320 6.800 656.040 1562.640 ;
    RECT 658.760 6.800 661.480 1562.640 ;
    RECT 664.200 6.800 666.920 1562.640 ;
    RECT 669.640 6.800 672.360 1562.640 ;
    RECT 675.080 6.800 677.800 1562.640 ;
    RECT 680.520 6.800 683.240 1562.640 ;
    RECT 685.960 6.800 688.680 1562.640 ;
    RECT 691.400 6.800 694.120 1562.640 ;
    RECT 696.840 6.800 699.560 1562.640 ;
    RECT 702.280 6.800 705.000 1562.640 ;
    RECT 707.720 6.800 710.440 1562.640 ;
    RECT 713.160 6.800 715.880 1562.640 ;
    RECT 718.600 6.800 721.320 1562.640 ;
    RECT 724.040 6.800 726.760 1562.640 ;
    RECT 729.480 6.800 732.200 1562.640 ;
    RECT 734.920 6.800 737.640 1562.640 ;
    RECT 740.360 6.800 743.080 1562.640 ;
    RECT 745.800 6.800 748.520 1562.640 ;
    RECT 751.240 6.800 753.960 1562.640 ;
    RECT 756.680 6.800 759.400 1562.640 ;
    RECT 762.120 6.800 764.840 1562.640 ;
    RECT 767.560 6.800 770.280 1562.640 ;
    RECT 773.000 6.800 775.720 1562.640 ;
    RECT 778.440 6.800 781.160 1562.640 ;
    RECT 783.880 6.800 786.600 1562.640 ;
    RECT 789.320 6.800 792.040 1562.640 ;
    RECT 794.760 6.800 797.480 1562.640 ;
    RECT 800.200 6.800 802.920 1562.640 ;
    RECT 805.640 6.800 808.360 1562.640 ;
    RECT 811.080 6.800 813.800 1562.640 ;
    RECT 816.520 6.800 819.240 1562.640 ;
    RECT 821.960 6.800 824.680 1562.640 ;
    RECT 827.400 6.800 830.120 1562.640 ;
    RECT 832.840 6.800 835.560 1562.640 ;
    RECT 838.280 6.800 841.000 1562.640 ;
    RECT 843.720 6.800 846.440 1562.640 ;
    RECT 849.160 6.800 851.880 1562.640 ;
    RECT 854.600 6.800 857.320 1562.640 ;
    RECT 860.040 6.800 862.760 1562.640 ;
    RECT 865.480 6.800 868.200 1562.640 ;
    RECT 870.920 6.800 873.640 1562.640 ;
    RECT 876.360 6.800 879.080 1562.640 ;
    RECT 881.800 6.800 884.520 1562.640 ;
    RECT 887.240 6.800 889.960 1562.640 ;
    RECT 892.680 6.800 895.400 1562.640 ;
    RECT 898.120 6.800 900.840 1562.640 ;
    RECT 903.560 6.800 906.280 1562.640 ;
    RECT 909.000 6.800 911.720 1562.640 ;
    RECT 914.440 6.800 917.160 1562.640 ;
    RECT 919.880 6.800 922.600 1562.640 ;
    RECT 925.320 6.800 928.040 1562.640 ;
    RECT 930.760 6.800 933.480 1562.640 ;
    RECT 936.200 6.800 938.920 1562.640 ;
    RECT 941.640 6.800 944.360 1562.640 ;
    RECT 947.080 6.800 949.800 1562.640 ;
    RECT 952.520 6.800 955.240 1562.640 ;
    RECT 957.960 6.800 960.680 1562.640 ;
    RECT 963.400 6.800 966.120 1562.640 ;
    RECT 968.840 6.800 971.560 1562.640 ;
    RECT 974.280 6.800 977.000 1562.640 ;
    RECT 979.720 6.800 982.440 1562.640 ;
    RECT 985.160 6.800 987.880 1562.640 ;
    RECT 990.600 6.800 993.320 1562.640 ;
    RECT 996.040 6.800 998.760 1562.640 ;
    RECT 1001.480 6.800 1004.200 1562.640 ;
    RECT 1006.920 6.800 1009.640 1562.640 ;
    RECT 1012.360 6.800 1015.080 1562.640 ;
    RECT 1017.800 6.800 1020.520 1562.640 ;
    RECT 1023.240 6.800 1025.960 1562.640 ;
    RECT 1028.680 6.800 1031.400 1562.640 ;
    RECT 1034.120 6.800 1036.840 1562.640 ;
    RECT 1039.560 6.800 1042.280 1562.640 ;
    RECT 1045.000 6.800 1047.720 1562.640 ;
    RECT 1050.440 6.800 1053.160 1562.640 ;
    RECT 1055.880 6.800 1058.600 1562.640 ;
    RECT 1061.320 6.800 1064.040 1562.640 ;
    RECT 1066.760 6.800 1069.480 1562.640 ;
    RECT 1072.200 6.800 1074.920 1562.640 ;
    RECT 1077.640 6.800 1080.360 1562.640 ;
    RECT 1083.080 6.800 1085.800 1562.640 ;
    RECT 1088.520 6.800 1091.240 1562.640 ;
    RECT 1093.960 6.800 1096.680 1562.640 ;
    RECT 1099.400 6.800 1102.120 1562.640 ;
    RECT 1104.840 6.800 1107.560 1562.640 ;
    RECT 1110.280 6.800 1113.000 1562.640 ;
    RECT 1115.720 6.800 1118.440 1562.640 ;
    RECT 1121.160 6.800 1123.880 1562.640 ;
    RECT 1126.600 6.800 1129.320 1562.640 ;
    RECT 1132.040 6.800 1134.760 1562.640 ;
    RECT 1137.480 6.800 1140.200 1562.640 ;
    RECT 1142.920 6.800 1145.640 1562.640 ;
    RECT 1148.360 6.800 1151.080 1562.640 ;
    RECT 1153.800 6.800 1156.520 1562.640 ;
    RECT 1159.240 6.800 1161.960 1562.640 ;
    RECT 1164.680 6.800 1167.400 1562.640 ;
    RECT 1170.120 6.800 1172.840 1562.640 ;
    RECT 1175.560 6.800 1178.280 1562.640 ;
    RECT 1181.000 6.800 1183.720 1562.640 ;
    RECT 1186.440 6.800 1189.160 1562.640 ;
    RECT 1191.880 6.800 1194.600 1562.640 ;
    RECT 1197.320 6.800 1200.040 1562.640 ;
    RECT 1202.760 6.800 1205.480 1562.640 ;
    RECT 1208.200 6.800 1210.920 1562.640 ;
    RECT 1213.640 6.800 1216.360 1562.640 ;
    RECT 1219.080 6.800 1221.800 1562.640 ;
    RECT 1224.520 6.800 1227.240 1562.640 ;
    RECT 1229.960 6.800 1232.680 1562.640 ;
    RECT 1235.400 6.800 1238.120 1562.640 ;
    RECT 1240.840 6.800 1243.560 1562.640 ;
    RECT 1246.280 6.800 1249.000 1562.640 ;
    RECT 1251.720 6.800 1254.440 1562.640 ;
    RECT 1257.160 6.800 1259.880 1562.640 ;
    RECT 1262.600 6.800 1265.320 1562.640 ;
    RECT 1268.040 6.800 1270.760 1562.640 ;
    RECT 1273.480 6.800 1276.200 1562.640 ;
    RECT 1278.920 6.800 1281.640 1562.640 ;
    RECT 1284.360 6.800 1287.080 1562.640 ;
    RECT 1289.800 6.800 1292.520 1562.640 ;
    RECT 1295.240 6.800 1302.720 1562.640 ;
    LAYER OVERLAP ;
    RECT 0 0 1302.720 1569.440 ;
  END
END fakeram_512x256_1r1w

END LIBRARY
