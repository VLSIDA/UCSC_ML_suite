VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_1x256_1r1w
  FOREIGN sram_1x256_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 130.910 BY 163.800 ;
  CLASS BLOCK ;
  PIN w_mask_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 -10.115 0.070 -10.045 ;
    END
  END w_mask_w1[0]
  PIN rd_out_r1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 -10.115 0.070 -10.045 ;
    END
  END rd_out_r1[0]
  PIN wd_in_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 -10.115 0.070 -10.045 ;
    END
  END wd_in_w1[0]
  PIN addr_w1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 -10.115 0.070 -10.045 ;
    END
  END addr_w1[0]
  PIN addr_w1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END addr_w1[1]
  PIN addr_w1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.845 0.070 12.915 ;
    END
  END addr_w1[2]
  PIN addr_w1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END addr_w1[3]
  PIN addr_w1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.805 0.070 35.875 ;
    END
  END addr_w1[4]
  PIN addr_w1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.285 0.070 47.355 ;
    END
  END addr_w1[5]
  PIN addr_w1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END addr_w1[6]
  PIN addr_w1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.245 0.070 70.315 ;
    END
  END addr_w1[7]
  PIN addr_r1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.245 0.070 70.315 ;
    END
  END addr_r1[0]
  PIN addr_r1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.725 0.070 81.795 ;
    END
  END addr_r1[1]
  PIN addr_r1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.205 0.070 93.275 ;
    END
  END addr_r1[2]
  PIN addr_r1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.685 0.070 104.755 ;
    END
  END addr_r1[3]
  PIN addr_r1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.165 0.070 116.235 ;
    END
  END addr_r1[4]
  PIN addr_r1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.645 0.070 127.715 ;
    END
  END addr_r1[5]
  PIN addr_r1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.125 0.070 139.195 ;
    END
  END addr_r1[6]
  PIN addr_r1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.605 0.070 150.675 ;
    END
  END addr_r1[7]
  PIN we_in_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.605 0.070 150.675 ;
    END
  END we_in_w1
  PIN ce_w1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.125 0.070 139.195 ;
    END
  END ce_w1
  PIN ce_r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.125 0.070 139.195 ;
    END
  END ce_r1
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.125 0.070 139.195 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 162.400 ;
      RECT 3.500 1.400 3.780 162.400 ;
      RECT 5.740 1.400 6.020 162.400 ;
      RECT 7.980 1.400 8.260 162.400 ;
      RECT 10.220 1.400 10.500 162.400 ;
      RECT 12.460 1.400 12.740 162.400 ;
      RECT 14.700 1.400 14.980 162.400 ;
      RECT 16.940 1.400 17.220 162.400 ;
      RECT 19.180 1.400 19.460 162.400 ;
      RECT 21.420 1.400 21.700 162.400 ;
      RECT 23.660 1.400 23.940 162.400 ;
      RECT 25.900 1.400 26.180 162.400 ;
      RECT 28.140 1.400 28.420 162.400 ;
      RECT 30.380 1.400 30.660 162.400 ;
      RECT 32.620 1.400 32.900 162.400 ;
      RECT 34.860 1.400 35.140 162.400 ;
      RECT 37.100 1.400 37.380 162.400 ;
      RECT 39.340 1.400 39.620 162.400 ;
      RECT 41.580 1.400 41.860 162.400 ;
      RECT 43.820 1.400 44.100 162.400 ;
      RECT 46.060 1.400 46.340 162.400 ;
      RECT 48.300 1.400 48.580 162.400 ;
      RECT 50.540 1.400 50.820 162.400 ;
      RECT 52.780 1.400 53.060 162.400 ;
      RECT 55.020 1.400 55.300 162.400 ;
      RECT 57.260 1.400 57.540 162.400 ;
      RECT 59.500 1.400 59.780 162.400 ;
      RECT 61.740 1.400 62.020 162.400 ;
      RECT 63.980 1.400 64.260 162.400 ;
      RECT 66.220 1.400 66.500 162.400 ;
      RECT 68.460 1.400 68.740 162.400 ;
      RECT 70.700 1.400 70.980 162.400 ;
      RECT 72.940 1.400 73.220 162.400 ;
      RECT 75.180 1.400 75.460 162.400 ;
      RECT 77.420 1.400 77.700 162.400 ;
      RECT 79.660 1.400 79.940 162.400 ;
      RECT 81.900 1.400 82.180 162.400 ;
      RECT 84.140 1.400 84.420 162.400 ;
      RECT 86.380 1.400 86.660 162.400 ;
      RECT 88.620 1.400 88.900 162.400 ;
      RECT 90.860 1.400 91.140 162.400 ;
      RECT 93.100 1.400 93.380 162.400 ;
      RECT 95.340 1.400 95.620 162.400 ;
      RECT 97.580 1.400 97.860 162.400 ;
      RECT 99.820 1.400 100.100 162.400 ;
      RECT 102.060 1.400 102.340 162.400 ;
      RECT 104.300 1.400 104.580 162.400 ;
      RECT 106.540 1.400 106.820 162.400 ;
      RECT 108.780 1.400 109.060 162.400 ;
      RECT 111.020 1.400 111.300 162.400 ;
      RECT 113.260 1.400 113.540 162.400 ;
      RECT 115.500 1.400 115.780 162.400 ;
      RECT 117.740 1.400 118.020 162.400 ;
      RECT 119.980 1.400 120.260 162.400 ;
      RECT 122.220 1.400 122.500 162.400 ;
      RECT 124.460 1.400 124.740 162.400 ;
      RECT 126.700 1.400 126.980 162.400 ;
      RECT 128.940 1.400 129.220 162.400 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 162.400 ;
      RECT 4.620 1.400 4.900 162.400 ;
      RECT 6.860 1.400 7.140 162.400 ;
      RECT 9.100 1.400 9.380 162.400 ;
      RECT 11.340 1.400 11.620 162.400 ;
      RECT 13.580 1.400 13.860 162.400 ;
      RECT 15.820 1.400 16.100 162.400 ;
      RECT 18.060 1.400 18.340 162.400 ;
      RECT 20.300 1.400 20.580 162.400 ;
      RECT 22.540 1.400 22.820 162.400 ;
      RECT 24.780 1.400 25.060 162.400 ;
      RECT 27.020 1.400 27.300 162.400 ;
      RECT 29.260 1.400 29.540 162.400 ;
      RECT 31.500 1.400 31.780 162.400 ;
      RECT 33.740 1.400 34.020 162.400 ;
      RECT 35.980 1.400 36.260 162.400 ;
      RECT 38.220 1.400 38.500 162.400 ;
      RECT 40.460 1.400 40.740 162.400 ;
      RECT 42.700 1.400 42.980 162.400 ;
      RECT 44.940 1.400 45.220 162.400 ;
      RECT 47.180 1.400 47.460 162.400 ;
      RECT 49.420 1.400 49.700 162.400 ;
      RECT 51.660 1.400 51.940 162.400 ;
      RECT 53.900 1.400 54.180 162.400 ;
      RECT 56.140 1.400 56.420 162.400 ;
      RECT 58.380 1.400 58.660 162.400 ;
      RECT 60.620 1.400 60.900 162.400 ;
      RECT 62.860 1.400 63.140 162.400 ;
      RECT 65.100 1.400 65.380 162.400 ;
      RECT 67.340 1.400 67.620 162.400 ;
      RECT 69.580 1.400 69.860 162.400 ;
      RECT 71.820 1.400 72.100 162.400 ;
      RECT 74.060 1.400 74.340 162.400 ;
      RECT 76.300 1.400 76.580 162.400 ;
      RECT 78.540 1.400 78.820 162.400 ;
      RECT 80.780 1.400 81.060 162.400 ;
      RECT 83.020 1.400 83.300 162.400 ;
      RECT 85.260 1.400 85.540 162.400 ;
      RECT 87.500 1.400 87.780 162.400 ;
      RECT 89.740 1.400 90.020 162.400 ;
      RECT 91.980 1.400 92.260 162.400 ;
      RECT 94.220 1.400 94.500 162.400 ;
      RECT 96.460 1.400 96.740 162.400 ;
      RECT 98.700 1.400 98.980 162.400 ;
      RECT 100.940 1.400 101.220 162.400 ;
      RECT 103.180 1.400 103.460 162.400 ;
      RECT 105.420 1.400 105.700 162.400 ;
      RECT 107.660 1.400 107.940 162.400 ;
      RECT 109.900 1.400 110.180 162.400 ;
      RECT 112.140 1.400 112.420 162.400 ;
      RECT 114.380 1.400 114.660 162.400 ;
      RECT 116.620 1.400 116.900 162.400 ;
      RECT 118.860 1.400 119.140 162.400 ;
      RECT 121.100 1.400 121.380 162.400 ;
      RECT 123.340 1.400 123.620 162.400 ;
      RECT 125.580 1.400 125.860 162.400 ;
      RECT 127.820 1.400 128.100 162.400 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 130.910 163.800 ;
    LAYER metal2 ;
    RECT 0 0 130.910 163.800 ;
    LAYER metal3 ;
    RECT 0.070 0 130.910 163.800 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.365 ;
    RECT 0 1.435 0.070 1.365 ;
    RECT 0 1.435 0.070 1.365 ;
    RECT 0 1.435 0.070 12.845 ;
    RECT 0 12.915 0.070 24.325 ;
    RECT 0 24.395 0.070 35.805 ;
    RECT 0 35.875 0.070 47.285 ;
    RECT 0 47.355 0.070 58.765 ;
    RECT 0 58.835 0.070 70.245 ;
    RECT 0 70.315 0.070 81.725 ;
    RECT 0 81.795 0.070 81.725 ;
    RECT 0 81.795 0.070 93.205 ;
    RECT 0 93.275 0.070 104.685 ;
    RECT 0 104.755 0.070 163.800 ;
    LAYER metal4 ;
    RECT 0 0 130.910 1.400 ;
    RECT 0 162.400 130.910 163.800 ;
    RECT 0.000 1.400 1.260 162.400 ;
    RECT 1.540 1.400 2.380 162.400 ;
    RECT 2.660 1.400 3.500 162.400 ;
    RECT 3.780 1.400 4.620 162.400 ;
    RECT 4.900 1.400 5.740 162.400 ;
    RECT 6.020 1.400 6.860 162.400 ;
    RECT 7.140 1.400 7.980 162.400 ;
    RECT 8.260 1.400 9.100 162.400 ;
    RECT 9.380 1.400 10.220 162.400 ;
    RECT 10.500 1.400 11.340 162.400 ;
    RECT 11.620 1.400 12.460 162.400 ;
    RECT 12.740 1.400 13.580 162.400 ;
    RECT 13.860 1.400 14.700 162.400 ;
    RECT 14.980 1.400 15.820 162.400 ;
    RECT 16.100 1.400 16.940 162.400 ;
    RECT 17.220 1.400 18.060 162.400 ;
    RECT 18.340 1.400 19.180 162.400 ;
    RECT 19.460 1.400 20.300 162.400 ;
    RECT 20.580 1.400 21.420 162.400 ;
    RECT 21.700 1.400 22.540 162.400 ;
    RECT 22.820 1.400 23.660 162.400 ;
    RECT 23.940 1.400 24.780 162.400 ;
    RECT 25.060 1.400 25.900 162.400 ;
    RECT 26.180 1.400 27.020 162.400 ;
    RECT 27.300 1.400 28.140 162.400 ;
    RECT 28.420 1.400 29.260 162.400 ;
    RECT 29.540 1.400 30.380 162.400 ;
    RECT 30.660 1.400 31.500 162.400 ;
    RECT 31.780 1.400 32.620 162.400 ;
    RECT 32.900 1.400 33.740 162.400 ;
    RECT 34.020 1.400 34.860 162.400 ;
    RECT 35.140 1.400 35.980 162.400 ;
    RECT 36.260 1.400 37.100 162.400 ;
    RECT 37.380 1.400 38.220 162.400 ;
    RECT 38.500 1.400 39.340 162.400 ;
    RECT 39.620 1.400 40.460 162.400 ;
    RECT 40.740 1.400 41.580 162.400 ;
    RECT 41.860 1.400 42.700 162.400 ;
    RECT 42.980 1.400 43.820 162.400 ;
    RECT 44.100 1.400 44.940 162.400 ;
    RECT 45.220 1.400 46.060 162.400 ;
    RECT 46.340 1.400 47.180 162.400 ;
    RECT 47.460 1.400 48.300 162.400 ;
    RECT 48.580 1.400 49.420 162.400 ;
    RECT 49.700 1.400 50.540 162.400 ;
    RECT 50.820 1.400 51.660 162.400 ;
    RECT 51.940 1.400 52.780 162.400 ;
    RECT 53.060 1.400 53.900 162.400 ;
    RECT 54.180 1.400 55.020 162.400 ;
    RECT 55.300 1.400 56.140 162.400 ;
    RECT 56.420 1.400 57.260 162.400 ;
    RECT 57.540 1.400 58.380 162.400 ;
    RECT 58.660 1.400 59.500 162.400 ;
    RECT 59.780 1.400 60.620 162.400 ;
    RECT 60.900 1.400 61.740 162.400 ;
    RECT 62.020 1.400 62.860 162.400 ;
    RECT 63.140 1.400 63.980 162.400 ;
    RECT 64.260 1.400 65.100 162.400 ;
    RECT 65.380 1.400 66.220 162.400 ;
    RECT 66.500 1.400 67.340 162.400 ;
    RECT 67.620 1.400 68.460 162.400 ;
    RECT 68.740 1.400 69.580 162.400 ;
    RECT 69.860 1.400 70.700 162.400 ;
    RECT 70.980 1.400 71.820 162.400 ;
    RECT 72.100 1.400 72.940 162.400 ;
    RECT 73.220 1.400 74.060 162.400 ;
    RECT 74.340 1.400 75.180 162.400 ;
    RECT 75.460 1.400 76.300 162.400 ;
    RECT 76.580 1.400 77.420 162.400 ;
    RECT 77.700 1.400 78.540 162.400 ;
    RECT 78.820 1.400 79.660 162.400 ;
    RECT 79.940 1.400 80.780 162.400 ;
    RECT 81.060 1.400 81.900 162.400 ;
    RECT 82.180 1.400 83.020 162.400 ;
    RECT 83.300 1.400 84.140 162.400 ;
    RECT 84.420 1.400 85.260 162.400 ;
    RECT 85.540 1.400 86.380 162.400 ;
    RECT 86.660 1.400 87.500 162.400 ;
    RECT 87.780 1.400 88.620 162.400 ;
    RECT 88.900 1.400 89.740 162.400 ;
    RECT 90.020 1.400 90.860 162.400 ;
    RECT 91.140 1.400 91.980 162.400 ;
    RECT 92.260 1.400 93.100 162.400 ;
    RECT 93.380 1.400 94.220 162.400 ;
    RECT 94.500 1.400 95.340 162.400 ;
    RECT 95.620 1.400 96.460 162.400 ;
    RECT 96.740 1.400 97.580 162.400 ;
    RECT 97.860 1.400 98.700 162.400 ;
    RECT 98.980 1.400 99.820 162.400 ;
    RECT 100.100 1.400 100.940 162.400 ;
    RECT 101.220 1.400 102.060 162.400 ;
    RECT 102.340 1.400 103.180 162.400 ;
    RECT 103.460 1.400 104.300 162.400 ;
    RECT 104.580 1.400 105.420 162.400 ;
    RECT 105.700 1.400 106.540 162.400 ;
    RECT 106.820 1.400 107.660 162.400 ;
    RECT 107.940 1.400 108.780 162.400 ;
    RECT 109.060 1.400 109.900 162.400 ;
    RECT 110.180 1.400 111.020 162.400 ;
    RECT 111.300 1.400 112.140 162.400 ;
    RECT 112.420 1.400 113.260 162.400 ;
    RECT 113.540 1.400 114.380 162.400 ;
    RECT 114.660 1.400 115.500 162.400 ;
    RECT 115.780 1.400 116.620 162.400 ;
    RECT 116.900 1.400 117.740 162.400 ;
    RECT 118.020 1.400 118.860 162.400 ;
    RECT 119.140 1.400 119.980 162.400 ;
    RECT 120.260 1.400 121.100 162.400 ;
    RECT 121.380 1.400 122.220 162.400 ;
    RECT 122.500 1.400 123.340 162.400 ;
    RECT 123.620 1.400 124.460 162.400 ;
    RECT 124.740 1.400 125.580 162.400 ;
    RECT 125.860 1.400 126.700 162.400 ;
    RECT 126.980 1.400 127.820 162.400 ;
    RECT 128.100 1.400 128.940 162.400 ;
    RECT 129.220 1.400 130.910 162.400 ;
    LAYER OVERLAP ;
    RECT 0 0 130.910 163.800 ;
  END
END sram_1x256_1r1w

END LIBRARY
