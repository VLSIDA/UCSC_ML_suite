VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_512x2048_1r1w
  FOREIGN fakeram_512x2048_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 1609.300 BY 1512.000 ;
  CLASS BLOCK ;
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 0.805 0.140 0.875 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.585 0.140 11.655 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.365 0.140 22.435 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.145 0.140 33.215 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.925 0.140 43.995 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.705 0.140 54.775 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.485 0.140 65.555 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.265 0.140 76.335 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.045 0.140 87.115 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.825 0.140 97.895 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.605 0.140 108.675 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.385 0.140 119.455 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.165 0.140 130.235 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.945 0.140 141.015 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.725 0.140 151.795 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.505 0.140 162.575 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.285 0.140 173.355 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.065 0.140 184.135 ;
    END
  END w0_wd_in[17]
  PIN w0_wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.845 0.140 194.915 ;
    END
  END w0_wd_in[18]
  PIN w0_wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.625 0.140 205.695 ;
    END
  END w0_wd_in[19]
  PIN w0_wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.405 0.140 216.475 ;
    END
  END w0_wd_in[20]
  PIN w0_wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.185 0.140 227.255 ;
    END
  END w0_wd_in[21]
  PIN w0_wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.965 0.140 238.035 ;
    END
  END w0_wd_in[22]
  PIN w0_wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.745 0.140 248.815 ;
    END
  END w0_wd_in[23]
  PIN w0_wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.525 0.140 259.595 ;
    END
  END w0_wd_in[24]
  PIN w0_wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.305 0.140 270.375 ;
    END
  END w0_wd_in[25]
  PIN w0_wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.085 0.140 281.155 ;
    END
  END w0_wd_in[26]
  PIN w0_wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.865 0.140 291.935 ;
    END
  END w0_wd_in[27]
  PIN w0_wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.645 0.140 302.715 ;
    END
  END w0_wd_in[28]
  PIN w0_wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.425 0.140 313.495 ;
    END
  END w0_wd_in[29]
  PIN w0_wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.205 0.140 324.275 ;
    END
  END w0_wd_in[30]
  PIN w0_wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.985 0.140 335.055 ;
    END
  END w0_wd_in[31]
  PIN w0_wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.765 0.140 345.835 ;
    END
  END w0_wd_in[32]
  PIN w0_wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.545 0.140 356.615 ;
    END
  END w0_wd_in[33]
  PIN w0_wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.325 0.140 367.395 ;
    END
  END w0_wd_in[34]
  PIN w0_wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.105 0.140 378.175 ;
    END
  END w0_wd_in[35]
  PIN w0_wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.885 0.140 388.955 ;
    END
  END w0_wd_in[36]
  PIN w0_wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.665 0.140 399.735 ;
    END
  END w0_wd_in[37]
  PIN w0_wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 410.445 0.140 410.515 ;
    END
  END w0_wd_in[38]
  PIN w0_wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 421.225 0.140 421.295 ;
    END
  END w0_wd_in[39]
  PIN w0_wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 432.005 0.140 432.075 ;
    END
  END w0_wd_in[40]
  PIN w0_wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 442.785 0.140 442.855 ;
    END
  END w0_wd_in[41]
  PIN w0_wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 453.565 0.140 453.635 ;
    END
  END w0_wd_in[42]
  PIN w0_wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 464.345 0.140 464.415 ;
    END
  END w0_wd_in[43]
  PIN w0_wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 475.125 0.140 475.195 ;
    END
  END w0_wd_in[44]
  PIN w0_wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 485.905 0.140 485.975 ;
    END
  END w0_wd_in[45]
  PIN w0_wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 496.685 0.140 496.755 ;
    END
  END w0_wd_in[46]
  PIN w0_wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.465 0.140 507.535 ;
    END
  END w0_wd_in[47]
  PIN w0_wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.245 0.140 518.315 ;
    END
  END w0_wd_in[48]
  PIN w0_wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.025 0.140 529.095 ;
    END
  END w0_wd_in[49]
  PIN w0_wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.805 0.140 539.875 ;
    END
  END w0_wd_in[50]
  PIN w0_wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.585 0.140 550.655 ;
    END
  END w0_wd_in[51]
  PIN w0_wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.365 0.140 561.435 ;
    END
  END w0_wd_in[52]
  PIN w0_wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.145 0.140 572.215 ;
    END
  END w0_wd_in[53]
  PIN w0_wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.925 0.140 582.995 ;
    END
  END w0_wd_in[54]
  PIN w0_wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.705 0.140 593.775 ;
    END
  END w0_wd_in[55]
  PIN w0_wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.485 0.140 604.555 ;
    END
  END w0_wd_in[56]
  PIN w0_wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.265 0.140 615.335 ;
    END
  END w0_wd_in[57]
  PIN w0_wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.045 0.140 626.115 ;
    END
  END w0_wd_in[58]
  PIN w0_wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.825 0.140 636.895 ;
    END
  END w0_wd_in[59]
  PIN w0_wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.605 0.140 647.675 ;
    END
  END w0_wd_in[60]
  PIN w0_wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.385 0.140 658.455 ;
    END
  END w0_wd_in[61]
  PIN w0_wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.165 0.140 669.235 ;
    END
  END w0_wd_in[62]
  PIN w0_wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.945 0.140 680.015 ;
    END
  END w0_wd_in[63]
  PIN w0_wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 690.725 0.140 690.795 ;
    END
  END w0_wd_in[64]
  PIN w0_wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.505 0.140 701.575 ;
    END
  END w0_wd_in[65]
  PIN w0_wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.285 0.140 712.355 ;
    END
  END w0_wd_in[66]
  PIN w0_wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.065 0.140 723.135 ;
    END
  END w0_wd_in[67]
  PIN w0_wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.845 0.140 733.915 ;
    END
  END w0_wd_in[68]
  PIN w0_wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 744.625 0.140 744.695 ;
    END
  END w0_wd_in[69]
  PIN w0_wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 755.405 0.140 755.475 ;
    END
  END w0_wd_in[70]
  PIN w0_wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 766.185 0.140 766.255 ;
    END
  END w0_wd_in[71]
  PIN w0_wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 776.965 0.140 777.035 ;
    END
  END w0_wd_in[72]
  PIN w0_wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 787.745 0.140 787.815 ;
    END
  END w0_wd_in[73]
  PIN w0_wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 798.525 0.140 798.595 ;
    END
  END w0_wd_in[74]
  PIN w0_wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 809.305 0.140 809.375 ;
    END
  END w0_wd_in[75]
  PIN w0_wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 820.085 0.140 820.155 ;
    END
  END w0_wd_in[76]
  PIN w0_wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 830.865 0.140 830.935 ;
    END
  END w0_wd_in[77]
  PIN w0_wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 841.645 0.140 841.715 ;
    END
  END w0_wd_in[78]
  PIN w0_wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.425 0.140 852.495 ;
    END
  END w0_wd_in[79]
  PIN w0_wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 863.205 0.140 863.275 ;
    END
  END w0_wd_in[80]
  PIN w0_wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.985 0.140 874.055 ;
    END
  END w0_wd_in[81]
  PIN w0_wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 884.765 0.140 884.835 ;
    END
  END w0_wd_in[82]
  PIN w0_wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 895.545 0.140 895.615 ;
    END
  END w0_wd_in[83]
  PIN w0_wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 906.325 0.140 906.395 ;
    END
  END w0_wd_in[84]
  PIN w0_wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 917.105 0.140 917.175 ;
    END
  END w0_wd_in[85]
  PIN w0_wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 927.885 0.140 927.955 ;
    END
  END w0_wd_in[86]
  PIN w0_wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 938.665 0.140 938.735 ;
    END
  END w0_wd_in[87]
  PIN w0_wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 949.445 0.140 949.515 ;
    END
  END w0_wd_in[88]
  PIN w0_wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 960.225 0.140 960.295 ;
    END
  END w0_wd_in[89]
  PIN w0_wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 971.005 0.140 971.075 ;
    END
  END w0_wd_in[90]
  PIN w0_wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 981.785 0.140 981.855 ;
    END
  END w0_wd_in[91]
  PIN w0_wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 992.565 0.140 992.635 ;
    END
  END w0_wd_in[92]
  PIN w0_wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1003.345 0.140 1003.415 ;
    END
  END w0_wd_in[93]
  PIN w0_wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1014.125 0.140 1014.195 ;
    END
  END w0_wd_in[94]
  PIN w0_wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1024.905 0.140 1024.975 ;
    END
  END w0_wd_in[95]
  PIN w0_wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1035.685 0.140 1035.755 ;
    END
  END w0_wd_in[96]
  PIN w0_wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1046.465 0.140 1046.535 ;
    END
  END w0_wd_in[97]
  PIN w0_wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1057.245 0.140 1057.315 ;
    END
  END w0_wd_in[98]
  PIN w0_wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1068.025 0.140 1068.095 ;
    END
  END w0_wd_in[99]
  PIN w0_wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1078.805 0.140 1078.875 ;
    END
  END w0_wd_in[100]
  PIN w0_wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1089.585 0.140 1089.655 ;
    END
  END w0_wd_in[101]
  PIN w0_wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1100.365 0.140 1100.435 ;
    END
  END w0_wd_in[102]
  PIN w0_wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1111.145 0.140 1111.215 ;
    END
  END w0_wd_in[103]
  PIN w0_wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1121.925 0.140 1121.995 ;
    END
  END w0_wd_in[104]
  PIN w0_wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1132.705 0.140 1132.775 ;
    END
  END w0_wd_in[105]
  PIN w0_wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1143.485 0.140 1143.555 ;
    END
  END w0_wd_in[106]
  PIN w0_wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1154.265 0.140 1154.335 ;
    END
  END w0_wd_in[107]
  PIN w0_wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1165.045 0.140 1165.115 ;
    END
  END w0_wd_in[108]
  PIN w0_wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1175.825 0.140 1175.895 ;
    END
  END w0_wd_in[109]
  PIN w0_wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1186.605 0.140 1186.675 ;
    END
  END w0_wd_in[110]
  PIN w0_wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1197.385 0.140 1197.455 ;
    END
  END w0_wd_in[111]
  PIN w0_wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1208.165 0.140 1208.235 ;
    END
  END w0_wd_in[112]
  PIN w0_wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1218.945 0.140 1219.015 ;
    END
  END w0_wd_in[113]
  PIN w0_wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1229.725 0.140 1229.795 ;
    END
  END w0_wd_in[114]
  PIN w0_wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1240.505 0.140 1240.575 ;
    END
  END w0_wd_in[115]
  PIN w0_wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1251.285 0.140 1251.355 ;
    END
  END w0_wd_in[116]
  PIN w0_wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1262.065 0.140 1262.135 ;
    END
  END w0_wd_in[117]
  PIN w0_wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1272.845 0.140 1272.915 ;
    END
  END w0_wd_in[118]
  PIN w0_wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1283.625 0.140 1283.695 ;
    END
  END w0_wd_in[119]
  PIN w0_wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1294.405 0.140 1294.475 ;
    END
  END w0_wd_in[120]
  PIN w0_wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1305.185 0.140 1305.255 ;
    END
  END w0_wd_in[121]
  PIN w0_wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1315.965 0.140 1316.035 ;
    END
  END w0_wd_in[122]
  PIN w0_wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1326.745 0.140 1326.815 ;
    END
  END w0_wd_in[123]
  PIN w0_wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1337.525 0.140 1337.595 ;
    END
  END w0_wd_in[124]
  PIN w0_wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1348.305 0.140 1348.375 ;
    END
  END w0_wd_in[125]
  PIN w0_wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1359.085 0.140 1359.155 ;
    END
  END w0_wd_in[126]
  PIN w0_wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1369.865 0.140 1369.935 ;
    END
  END w0_wd_in[127]
  PIN w0_wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 0.805 1609.300 0.875 ;
    END
  END w0_wd_in[128]
  PIN w0_wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 11.585 1609.300 11.655 ;
    END
  END w0_wd_in[129]
  PIN w0_wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 22.365 1609.300 22.435 ;
    END
  END w0_wd_in[130]
  PIN w0_wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 33.145 1609.300 33.215 ;
    END
  END w0_wd_in[131]
  PIN w0_wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 43.925 1609.300 43.995 ;
    END
  END w0_wd_in[132]
  PIN w0_wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 54.705 1609.300 54.775 ;
    END
  END w0_wd_in[133]
  PIN w0_wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 65.485 1609.300 65.555 ;
    END
  END w0_wd_in[134]
  PIN w0_wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 76.265 1609.300 76.335 ;
    END
  END w0_wd_in[135]
  PIN w0_wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 87.045 1609.300 87.115 ;
    END
  END w0_wd_in[136]
  PIN w0_wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 97.825 1609.300 97.895 ;
    END
  END w0_wd_in[137]
  PIN w0_wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 108.605 1609.300 108.675 ;
    END
  END w0_wd_in[138]
  PIN w0_wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 119.385 1609.300 119.455 ;
    END
  END w0_wd_in[139]
  PIN w0_wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 130.165 1609.300 130.235 ;
    END
  END w0_wd_in[140]
  PIN w0_wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 140.945 1609.300 141.015 ;
    END
  END w0_wd_in[141]
  PIN w0_wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 151.725 1609.300 151.795 ;
    END
  END w0_wd_in[142]
  PIN w0_wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 162.505 1609.300 162.575 ;
    END
  END w0_wd_in[143]
  PIN w0_wd_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 173.285 1609.300 173.355 ;
    END
  END w0_wd_in[144]
  PIN w0_wd_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 184.065 1609.300 184.135 ;
    END
  END w0_wd_in[145]
  PIN w0_wd_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 194.845 1609.300 194.915 ;
    END
  END w0_wd_in[146]
  PIN w0_wd_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 205.625 1609.300 205.695 ;
    END
  END w0_wd_in[147]
  PIN w0_wd_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 216.405 1609.300 216.475 ;
    END
  END w0_wd_in[148]
  PIN w0_wd_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 227.185 1609.300 227.255 ;
    END
  END w0_wd_in[149]
  PIN w0_wd_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 237.965 1609.300 238.035 ;
    END
  END w0_wd_in[150]
  PIN w0_wd_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 248.745 1609.300 248.815 ;
    END
  END w0_wd_in[151]
  PIN w0_wd_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 259.525 1609.300 259.595 ;
    END
  END w0_wd_in[152]
  PIN w0_wd_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 270.305 1609.300 270.375 ;
    END
  END w0_wd_in[153]
  PIN w0_wd_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 281.085 1609.300 281.155 ;
    END
  END w0_wd_in[154]
  PIN w0_wd_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 291.865 1609.300 291.935 ;
    END
  END w0_wd_in[155]
  PIN w0_wd_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 302.645 1609.300 302.715 ;
    END
  END w0_wd_in[156]
  PIN w0_wd_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 313.425 1609.300 313.495 ;
    END
  END w0_wd_in[157]
  PIN w0_wd_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 324.205 1609.300 324.275 ;
    END
  END w0_wd_in[158]
  PIN w0_wd_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 334.985 1609.300 335.055 ;
    END
  END w0_wd_in[159]
  PIN w0_wd_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 345.765 1609.300 345.835 ;
    END
  END w0_wd_in[160]
  PIN w0_wd_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 356.545 1609.300 356.615 ;
    END
  END w0_wd_in[161]
  PIN w0_wd_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 367.325 1609.300 367.395 ;
    END
  END w0_wd_in[162]
  PIN w0_wd_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 378.105 1609.300 378.175 ;
    END
  END w0_wd_in[163]
  PIN w0_wd_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 388.885 1609.300 388.955 ;
    END
  END w0_wd_in[164]
  PIN w0_wd_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 399.665 1609.300 399.735 ;
    END
  END w0_wd_in[165]
  PIN w0_wd_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 410.445 1609.300 410.515 ;
    END
  END w0_wd_in[166]
  PIN w0_wd_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 421.225 1609.300 421.295 ;
    END
  END w0_wd_in[167]
  PIN w0_wd_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 432.005 1609.300 432.075 ;
    END
  END w0_wd_in[168]
  PIN w0_wd_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 442.785 1609.300 442.855 ;
    END
  END w0_wd_in[169]
  PIN w0_wd_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 453.565 1609.300 453.635 ;
    END
  END w0_wd_in[170]
  PIN w0_wd_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 464.345 1609.300 464.415 ;
    END
  END w0_wd_in[171]
  PIN w0_wd_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 475.125 1609.300 475.195 ;
    END
  END w0_wd_in[172]
  PIN w0_wd_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 485.905 1609.300 485.975 ;
    END
  END w0_wd_in[173]
  PIN w0_wd_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 496.685 1609.300 496.755 ;
    END
  END w0_wd_in[174]
  PIN w0_wd_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 507.465 1609.300 507.535 ;
    END
  END w0_wd_in[175]
  PIN w0_wd_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 518.245 1609.300 518.315 ;
    END
  END w0_wd_in[176]
  PIN w0_wd_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 529.025 1609.300 529.095 ;
    END
  END w0_wd_in[177]
  PIN w0_wd_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 539.805 1609.300 539.875 ;
    END
  END w0_wd_in[178]
  PIN w0_wd_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 550.585 1609.300 550.655 ;
    END
  END w0_wd_in[179]
  PIN w0_wd_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 561.365 1609.300 561.435 ;
    END
  END w0_wd_in[180]
  PIN w0_wd_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 572.145 1609.300 572.215 ;
    END
  END w0_wd_in[181]
  PIN w0_wd_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 582.925 1609.300 582.995 ;
    END
  END w0_wd_in[182]
  PIN w0_wd_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 593.705 1609.300 593.775 ;
    END
  END w0_wd_in[183]
  PIN w0_wd_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 604.485 1609.300 604.555 ;
    END
  END w0_wd_in[184]
  PIN w0_wd_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 615.265 1609.300 615.335 ;
    END
  END w0_wd_in[185]
  PIN w0_wd_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 626.045 1609.300 626.115 ;
    END
  END w0_wd_in[186]
  PIN w0_wd_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 636.825 1609.300 636.895 ;
    END
  END w0_wd_in[187]
  PIN w0_wd_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 647.605 1609.300 647.675 ;
    END
  END w0_wd_in[188]
  PIN w0_wd_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 658.385 1609.300 658.455 ;
    END
  END w0_wd_in[189]
  PIN w0_wd_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 669.165 1609.300 669.235 ;
    END
  END w0_wd_in[190]
  PIN w0_wd_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 679.945 1609.300 680.015 ;
    END
  END w0_wd_in[191]
  PIN w0_wd_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 690.725 1609.300 690.795 ;
    END
  END w0_wd_in[192]
  PIN w0_wd_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 701.505 1609.300 701.575 ;
    END
  END w0_wd_in[193]
  PIN w0_wd_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 712.285 1609.300 712.355 ;
    END
  END w0_wd_in[194]
  PIN w0_wd_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 723.065 1609.300 723.135 ;
    END
  END w0_wd_in[195]
  PIN w0_wd_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 733.845 1609.300 733.915 ;
    END
  END w0_wd_in[196]
  PIN w0_wd_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 744.625 1609.300 744.695 ;
    END
  END w0_wd_in[197]
  PIN w0_wd_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 755.405 1609.300 755.475 ;
    END
  END w0_wd_in[198]
  PIN w0_wd_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 766.185 1609.300 766.255 ;
    END
  END w0_wd_in[199]
  PIN w0_wd_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 776.965 1609.300 777.035 ;
    END
  END w0_wd_in[200]
  PIN w0_wd_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 787.745 1609.300 787.815 ;
    END
  END w0_wd_in[201]
  PIN w0_wd_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 798.525 1609.300 798.595 ;
    END
  END w0_wd_in[202]
  PIN w0_wd_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 809.305 1609.300 809.375 ;
    END
  END w0_wd_in[203]
  PIN w0_wd_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 820.085 1609.300 820.155 ;
    END
  END w0_wd_in[204]
  PIN w0_wd_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 830.865 1609.300 830.935 ;
    END
  END w0_wd_in[205]
  PIN w0_wd_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 841.645 1609.300 841.715 ;
    END
  END w0_wd_in[206]
  PIN w0_wd_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 852.425 1609.300 852.495 ;
    END
  END w0_wd_in[207]
  PIN w0_wd_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 863.205 1609.300 863.275 ;
    END
  END w0_wd_in[208]
  PIN w0_wd_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 873.985 1609.300 874.055 ;
    END
  END w0_wd_in[209]
  PIN w0_wd_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 884.765 1609.300 884.835 ;
    END
  END w0_wd_in[210]
  PIN w0_wd_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 895.545 1609.300 895.615 ;
    END
  END w0_wd_in[211]
  PIN w0_wd_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 906.325 1609.300 906.395 ;
    END
  END w0_wd_in[212]
  PIN w0_wd_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 917.105 1609.300 917.175 ;
    END
  END w0_wd_in[213]
  PIN w0_wd_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 927.885 1609.300 927.955 ;
    END
  END w0_wd_in[214]
  PIN w0_wd_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 938.665 1609.300 938.735 ;
    END
  END w0_wd_in[215]
  PIN w0_wd_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 949.445 1609.300 949.515 ;
    END
  END w0_wd_in[216]
  PIN w0_wd_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 960.225 1609.300 960.295 ;
    END
  END w0_wd_in[217]
  PIN w0_wd_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 971.005 1609.300 971.075 ;
    END
  END w0_wd_in[218]
  PIN w0_wd_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 981.785 1609.300 981.855 ;
    END
  END w0_wd_in[219]
  PIN w0_wd_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 992.565 1609.300 992.635 ;
    END
  END w0_wd_in[220]
  PIN w0_wd_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1003.345 1609.300 1003.415 ;
    END
  END w0_wd_in[221]
  PIN w0_wd_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1014.125 1609.300 1014.195 ;
    END
  END w0_wd_in[222]
  PIN w0_wd_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1024.905 1609.300 1024.975 ;
    END
  END w0_wd_in[223]
  PIN w0_wd_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1035.685 1609.300 1035.755 ;
    END
  END w0_wd_in[224]
  PIN w0_wd_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1046.465 1609.300 1046.535 ;
    END
  END w0_wd_in[225]
  PIN w0_wd_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1057.245 1609.300 1057.315 ;
    END
  END w0_wd_in[226]
  PIN w0_wd_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1068.025 1609.300 1068.095 ;
    END
  END w0_wd_in[227]
  PIN w0_wd_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1078.805 1609.300 1078.875 ;
    END
  END w0_wd_in[228]
  PIN w0_wd_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1089.585 1609.300 1089.655 ;
    END
  END w0_wd_in[229]
  PIN w0_wd_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1100.365 1609.300 1100.435 ;
    END
  END w0_wd_in[230]
  PIN w0_wd_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1111.145 1609.300 1111.215 ;
    END
  END w0_wd_in[231]
  PIN w0_wd_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1121.925 1609.300 1121.995 ;
    END
  END w0_wd_in[232]
  PIN w0_wd_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1132.705 1609.300 1132.775 ;
    END
  END w0_wd_in[233]
  PIN w0_wd_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1143.485 1609.300 1143.555 ;
    END
  END w0_wd_in[234]
  PIN w0_wd_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1154.265 1609.300 1154.335 ;
    END
  END w0_wd_in[235]
  PIN w0_wd_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1165.045 1609.300 1165.115 ;
    END
  END w0_wd_in[236]
  PIN w0_wd_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1175.825 1609.300 1175.895 ;
    END
  END w0_wd_in[237]
  PIN w0_wd_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1186.605 1609.300 1186.675 ;
    END
  END w0_wd_in[238]
  PIN w0_wd_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1197.385 1609.300 1197.455 ;
    END
  END w0_wd_in[239]
  PIN w0_wd_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1208.165 1609.300 1208.235 ;
    END
  END w0_wd_in[240]
  PIN w0_wd_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1218.945 1609.300 1219.015 ;
    END
  END w0_wd_in[241]
  PIN w0_wd_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1229.725 1609.300 1229.795 ;
    END
  END w0_wd_in[242]
  PIN w0_wd_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1240.505 1609.300 1240.575 ;
    END
  END w0_wd_in[243]
  PIN w0_wd_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1251.285 1609.300 1251.355 ;
    END
  END w0_wd_in[244]
  PIN w0_wd_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1262.065 1609.300 1262.135 ;
    END
  END w0_wd_in[245]
  PIN w0_wd_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1272.845 1609.300 1272.915 ;
    END
  END w0_wd_in[246]
  PIN w0_wd_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1283.625 1609.300 1283.695 ;
    END
  END w0_wd_in[247]
  PIN w0_wd_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1294.405 1609.300 1294.475 ;
    END
  END w0_wd_in[248]
  PIN w0_wd_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1305.185 1609.300 1305.255 ;
    END
  END w0_wd_in[249]
  PIN w0_wd_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1315.965 1609.300 1316.035 ;
    END
  END w0_wd_in[250]
  PIN w0_wd_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1326.745 1609.300 1326.815 ;
    END
  END w0_wd_in[251]
  PIN w0_wd_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1337.525 1609.300 1337.595 ;
    END
  END w0_wd_in[252]
  PIN w0_wd_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1348.305 1609.300 1348.375 ;
    END
  END w0_wd_in[253]
  PIN w0_wd_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1359.085 1609.300 1359.155 ;
    END
  END w0_wd_in[254]
  PIN w0_wd_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1369.865 1609.300 1369.935 ;
    END
  END w0_wd_in[255]
  PIN w0_wd_in[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1.105 0.000 1.175 0.140 ;
    END
  END w0_wd_in[256]
  PIN w0_wd_in[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 4.145 0.000 4.215 0.140 ;
    END
  END w0_wd_in[257]
  PIN w0_wd_in[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 7.185 0.000 7.255 0.140 ;
    END
  END w0_wd_in[258]
  PIN w0_wd_in[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 10.225 0.000 10.295 0.140 ;
    END
  END w0_wd_in[259]
  PIN w0_wd_in[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 13.265 0.000 13.335 0.140 ;
    END
  END w0_wd_in[260]
  PIN w0_wd_in[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 16.305 0.000 16.375 0.140 ;
    END
  END w0_wd_in[261]
  PIN w0_wd_in[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 19.345 0.000 19.415 0.140 ;
    END
  END w0_wd_in[262]
  PIN w0_wd_in[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 22.385 0.000 22.455 0.140 ;
    END
  END w0_wd_in[263]
  PIN w0_wd_in[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 25.425 0.000 25.495 0.140 ;
    END
  END w0_wd_in[264]
  PIN w0_wd_in[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 28.465 0.000 28.535 0.140 ;
    END
  END w0_wd_in[265]
  PIN w0_wd_in[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 31.505 0.000 31.575 0.140 ;
    END
  END w0_wd_in[266]
  PIN w0_wd_in[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 34.545 0.000 34.615 0.140 ;
    END
  END w0_wd_in[267]
  PIN w0_wd_in[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 37.585 0.000 37.655 0.140 ;
    END
  END w0_wd_in[268]
  PIN w0_wd_in[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 40.625 0.000 40.695 0.140 ;
    END
  END w0_wd_in[269]
  PIN w0_wd_in[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 43.665 0.000 43.735 0.140 ;
    END
  END w0_wd_in[270]
  PIN w0_wd_in[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 46.705 0.000 46.775 0.140 ;
    END
  END w0_wd_in[271]
  PIN w0_wd_in[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 49.745 0.000 49.815 0.140 ;
    END
  END w0_wd_in[272]
  PIN w0_wd_in[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 52.785 0.000 52.855 0.140 ;
    END
  END w0_wd_in[273]
  PIN w0_wd_in[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 55.825 0.000 55.895 0.140 ;
    END
  END w0_wd_in[274]
  PIN w0_wd_in[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 58.865 0.000 58.935 0.140 ;
    END
  END w0_wd_in[275]
  PIN w0_wd_in[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 61.905 0.000 61.975 0.140 ;
    END
  END w0_wd_in[276]
  PIN w0_wd_in[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 64.945 0.000 65.015 0.140 ;
    END
  END w0_wd_in[277]
  PIN w0_wd_in[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 67.985 0.000 68.055 0.140 ;
    END
  END w0_wd_in[278]
  PIN w0_wd_in[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 71.025 0.000 71.095 0.140 ;
    END
  END w0_wd_in[279]
  PIN w0_wd_in[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 74.065 0.000 74.135 0.140 ;
    END
  END w0_wd_in[280]
  PIN w0_wd_in[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 77.105 0.000 77.175 0.140 ;
    END
  END w0_wd_in[281]
  PIN w0_wd_in[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 80.145 0.000 80.215 0.140 ;
    END
  END w0_wd_in[282]
  PIN w0_wd_in[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 83.185 0.000 83.255 0.140 ;
    END
  END w0_wd_in[283]
  PIN w0_wd_in[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 86.225 0.000 86.295 0.140 ;
    END
  END w0_wd_in[284]
  PIN w0_wd_in[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 89.265 0.000 89.335 0.140 ;
    END
  END w0_wd_in[285]
  PIN w0_wd_in[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 92.305 0.000 92.375 0.140 ;
    END
  END w0_wd_in[286]
  PIN w0_wd_in[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 95.345 0.000 95.415 0.140 ;
    END
  END w0_wd_in[287]
  PIN w0_wd_in[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 98.385 0.000 98.455 0.140 ;
    END
  END w0_wd_in[288]
  PIN w0_wd_in[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 101.425 0.000 101.495 0.140 ;
    END
  END w0_wd_in[289]
  PIN w0_wd_in[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 104.465 0.000 104.535 0.140 ;
    END
  END w0_wd_in[290]
  PIN w0_wd_in[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 107.505 0.000 107.575 0.140 ;
    END
  END w0_wd_in[291]
  PIN w0_wd_in[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 110.545 0.000 110.615 0.140 ;
    END
  END w0_wd_in[292]
  PIN w0_wd_in[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 113.585 0.000 113.655 0.140 ;
    END
  END w0_wd_in[293]
  PIN w0_wd_in[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 116.625 0.000 116.695 0.140 ;
    END
  END w0_wd_in[294]
  PIN w0_wd_in[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 119.665 0.000 119.735 0.140 ;
    END
  END w0_wd_in[295]
  PIN w0_wd_in[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 122.705 0.000 122.775 0.140 ;
    END
  END w0_wd_in[296]
  PIN w0_wd_in[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 125.745 0.000 125.815 0.140 ;
    END
  END w0_wd_in[297]
  PIN w0_wd_in[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 128.785 0.000 128.855 0.140 ;
    END
  END w0_wd_in[298]
  PIN w0_wd_in[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 131.825 0.000 131.895 0.140 ;
    END
  END w0_wd_in[299]
  PIN w0_wd_in[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 134.865 0.000 134.935 0.140 ;
    END
  END w0_wd_in[300]
  PIN w0_wd_in[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 137.905 0.000 137.975 0.140 ;
    END
  END w0_wd_in[301]
  PIN w0_wd_in[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 140.945 0.000 141.015 0.140 ;
    END
  END w0_wd_in[302]
  PIN w0_wd_in[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 143.985 0.000 144.055 0.140 ;
    END
  END w0_wd_in[303]
  PIN w0_wd_in[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 147.025 0.000 147.095 0.140 ;
    END
  END w0_wd_in[304]
  PIN w0_wd_in[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 150.065 0.000 150.135 0.140 ;
    END
  END w0_wd_in[305]
  PIN w0_wd_in[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 153.105 0.000 153.175 0.140 ;
    END
  END w0_wd_in[306]
  PIN w0_wd_in[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 156.145 0.000 156.215 0.140 ;
    END
  END w0_wd_in[307]
  PIN w0_wd_in[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 159.185 0.000 159.255 0.140 ;
    END
  END w0_wd_in[308]
  PIN w0_wd_in[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 162.225 0.000 162.295 0.140 ;
    END
  END w0_wd_in[309]
  PIN w0_wd_in[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 165.265 0.000 165.335 0.140 ;
    END
  END w0_wd_in[310]
  PIN w0_wd_in[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 168.305 0.000 168.375 0.140 ;
    END
  END w0_wd_in[311]
  PIN w0_wd_in[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 171.345 0.000 171.415 0.140 ;
    END
  END w0_wd_in[312]
  PIN w0_wd_in[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 174.385 0.000 174.455 0.140 ;
    END
  END w0_wd_in[313]
  PIN w0_wd_in[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 177.425 0.000 177.495 0.140 ;
    END
  END w0_wd_in[314]
  PIN w0_wd_in[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 180.465 0.000 180.535 0.140 ;
    END
  END w0_wd_in[315]
  PIN w0_wd_in[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 183.505 0.000 183.575 0.140 ;
    END
  END w0_wd_in[316]
  PIN w0_wd_in[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 186.545 0.000 186.615 0.140 ;
    END
  END w0_wd_in[317]
  PIN w0_wd_in[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 189.585 0.000 189.655 0.140 ;
    END
  END w0_wd_in[318]
  PIN w0_wd_in[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 192.625 0.000 192.695 0.140 ;
    END
  END w0_wd_in[319]
  PIN w0_wd_in[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 195.665 0.000 195.735 0.140 ;
    END
  END w0_wd_in[320]
  PIN w0_wd_in[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 198.705 0.000 198.775 0.140 ;
    END
  END w0_wd_in[321]
  PIN w0_wd_in[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 201.745 0.000 201.815 0.140 ;
    END
  END w0_wd_in[322]
  PIN w0_wd_in[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 204.785 0.000 204.855 0.140 ;
    END
  END w0_wd_in[323]
  PIN w0_wd_in[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 207.825 0.000 207.895 0.140 ;
    END
  END w0_wd_in[324]
  PIN w0_wd_in[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 210.865 0.000 210.935 0.140 ;
    END
  END w0_wd_in[325]
  PIN w0_wd_in[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 213.905 0.000 213.975 0.140 ;
    END
  END w0_wd_in[326]
  PIN w0_wd_in[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 216.945 0.000 217.015 0.140 ;
    END
  END w0_wd_in[327]
  PIN w0_wd_in[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 219.985 0.000 220.055 0.140 ;
    END
  END w0_wd_in[328]
  PIN w0_wd_in[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 223.025 0.000 223.095 0.140 ;
    END
  END w0_wd_in[329]
  PIN w0_wd_in[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 226.065 0.000 226.135 0.140 ;
    END
  END w0_wd_in[330]
  PIN w0_wd_in[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 229.105 0.000 229.175 0.140 ;
    END
  END w0_wd_in[331]
  PIN w0_wd_in[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 232.145 0.000 232.215 0.140 ;
    END
  END w0_wd_in[332]
  PIN w0_wd_in[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 235.185 0.000 235.255 0.140 ;
    END
  END w0_wd_in[333]
  PIN w0_wd_in[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 238.225 0.000 238.295 0.140 ;
    END
  END w0_wd_in[334]
  PIN w0_wd_in[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 241.265 0.000 241.335 0.140 ;
    END
  END w0_wd_in[335]
  PIN w0_wd_in[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 244.305 0.000 244.375 0.140 ;
    END
  END w0_wd_in[336]
  PIN w0_wd_in[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 247.345 0.000 247.415 0.140 ;
    END
  END w0_wd_in[337]
  PIN w0_wd_in[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 250.385 0.000 250.455 0.140 ;
    END
  END w0_wd_in[338]
  PIN w0_wd_in[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 253.425 0.000 253.495 0.140 ;
    END
  END w0_wd_in[339]
  PIN w0_wd_in[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 256.465 0.000 256.535 0.140 ;
    END
  END w0_wd_in[340]
  PIN w0_wd_in[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 259.505 0.000 259.575 0.140 ;
    END
  END w0_wd_in[341]
  PIN w0_wd_in[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 262.545 0.000 262.615 0.140 ;
    END
  END w0_wd_in[342]
  PIN w0_wd_in[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 265.585 0.000 265.655 0.140 ;
    END
  END w0_wd_in[343]
  PIN w0_wd_in[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 268.625 0.000 268.695 0.140 ;
    END
  END w0_wd_in[344]
  PIN w0_wd_in[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 271.665 0.000 271.735 0.140 ;
    END
  END w0_wd_in[345]
  PIN w0_wd_in[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 274.705 0.000 274.775 0.140 ;
    END
  END w0_wd_in[346]
  PIN w0_wd_in[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 277.745 0.000 277.815 0.140 ;
    END
  END w0_wd_in[347]
  PIN w0_wd_in[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 280.785 0.000 280.855 0.140 ;
    END
  END w0_wd_in[348]
  PIN w0_wd_in[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 283.825 0.000 283.895 0.140 ;
    END
  END w0_wd_in[349]
  PIN w0_wd_in[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 286.865 0.000 286.935 0.140 ;
    END
  END w0_wd_in[350]
  PIN w0_wd_in[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 289.905 0.000 289.975 0.140 ;
    END
  END w0_wd_in[351]
  PIN w0_wd_in[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 292.945 0.000 293.015 0.140 ;
    END
  END w0_wd_in[352]
  PIN w0_wd_in[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 295.985 0.000 296.055 0.140 ;
    END
  END w0_wd_in[353]
  PIN w0_wd_in[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 299.025 0.000 299.095 0.140 ;
    END
  END w0_wd_in[354]
  PIN w0_wd_in[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 302.065 0.000 302.135 0.140 ;
    END
  END w0_wd_in[355]
  PIN w0_wd_in[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 305.105 0.000 305.175 0.140 ;
    END
  END w0_wd_in[356]
  PIN w0_wd_in[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 308.145 0.000 308.215 0.140 ;
    END
  END w0_wd_in[357]
  PIN w0_wd_in[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 311.185 0.000 311.255 0.140 ;
    END
  END w0_wd_in[358]
  PIN w0_wd_in[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 314.225 0.000 314.295 0.140 ;
    END
  END w0_wd_in[359]
  PIN w0_wd_in[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 317.265 0.000 317.335 0.140 ;
    END
  END w0_wd_in[360]
  PIN w0_wd_in[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 320.305 0.000 320.375 0.140 ;
    END
  END w0_wd_in[361]
  PIN w0_wd_in[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 323.345 0.000 323.415 0.140 ;
    END
  END w0_wd_in[362]
  PIN w0_wd_in[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 326.385 0.000 326.455 0.140 ;
    END
  END w0_wd_in[363]
  PIN w0_wd_in[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 329.425 0.000 329.495 0.140 ;
    END
  END w0_wd_in[364]
  PIN w0_wd_in[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 332.465 0.000 332.535 0.140 ;
    END
  END w0_wd_in[365]
  PIN w0_wd_in[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 335.505 0.000 335.575 0.140 ;
    END
  END w0_wd_in[366]
  PIN w0_wd_in[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 338.545 0.000 338.615 0.140 ;
    END
  END w0_wd_in[367]
  PIN w0_wd_in[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 341.585 0.000 341.655 0.140 ;
    END
  END w0_wd_in[368]
  PIN w0_wd_in[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 344.625 0.000 344.695 0.140 ;
    END
  END w0_wd_in[369]
  PIN w0_wd_in[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 347.665 0.000 347.735 0.140 ;
    END
  END w0_wd_in[370]
  PIN w0_wd_in[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 350.705 0.000 350.775 0.140 ;
    END
  END w0_wd_in[371]
  PIN w0_wd_in[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 353.745 0.000 353.815 0.140 ;
    END
  END w0_wd_in[372]
  PIN w0_wd_in[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 356.785 0.000 356.855 0.140 ;
    END
  END w0_wd_in[373]
  PIN w0_wd_in[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 359.825 0.000 359.895 0.140 ;
    END
  END w0_wd_in[374]
  PIN w0_wd_in[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 362.865 0.000 362.935 0.140 ;
    END
  END w0_wd_in[375]
  PIN w0_wd_in[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 365.905 0.000 365.975 0.140 ;
    END
  END w0_wd_in[376]
  PIN w0_wd_in[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 368.945 0.000 369.015 0.140 ;
    END
  END w0_wd_in[377]
  PIN w0_wd_in[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 371.985 0.000 372.055 0.140 ;
    END
  END w0_wd_in[378]
  PIN w0_wd_in[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 375.025 0.000 375.095 0.140 ;
    END
  END w0_wd_in[379]
  PIN w0_wd_in[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 378.065 0.000 378.135 0.140 ;
    END
  END w0_wd_in[380]
  PIN w0_wd_in[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 381.105 0.000 381.175 0.140 ;
    END
  END w0_wd_in[381]
  PIN w0_wd_in[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 384.145 0.000 384.215 0.140 ;
    END
  END w0_wd_in[382]
  PIN w0_wd_in[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 387.185 0.000 387.255 0.140 ;
    END
  END w0_wd_in[383]
  PIN w0_wd_in[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 390.225 0.000 390.295 0.140 ;
    END
  END w0_wd_in[384]
  PIN w0_wd_in[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 393.265 0.000 393.335 0.140 ;
    END
  END w0_wd_in[385]
  PIN w0_wd_in[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 396.305 0.000 396.375 0.140 ;
    END
  END w0_wd_in[386]
  PIN w0_wd_in[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 399.345 0.000 399.415 0.140 ;
    END
  END w0_wd_in[387]
  PIN w0_wd_in[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 402.385 0.000 402.455 0.140 ;
    END
  END w0_wd_in[388]
  PIN w0_wd_in[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 405.425 0.000 405.495 0.140 ;
    END
  END w0_wd_in[389]
  PIN w0_wd_in[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 408.465 0.000 408.535 0.140 ;
    END
  END w0_wd_in[390]
  PIN w0_wd_in[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 411.505 0.000 411.575 0.140 ;
    END
  END w0_wd_in[391]
  PIN w0_wd_in[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 414.545 0.000 414.615 0.140 ;
    END
  END w0_wd_in[392]
  PIN w0_wd_in[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 417.585 0.000 417.655 0.140 ;
    END
  END w0_wd_in[393]
  PIN w0_wd_in[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 420.625 0.000 420.695 0.140 ;
    END
  END w0_wd_in[394]
  PIN w0_wd_in[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 423.665 0.000 423.735 0.140 ;
    END
  END w0_wd_in[395]
  PIN w0_wd_in[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 426.705 0.000 426.775 0.140 ;
    END
  END w0_wd_in[396]
  PIN w0_wd_in[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 429.745 0.000 429.815 0.140 ;
    END
  END w0_wd_in[397]
  PIN w0_wd_in[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 432.785 0.000 432.855 0.140 ;
    END
  END w0_wd_in[398]
  PIN w0_wd_in[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 435.825 0.000 435.895 0.140 ;
    END
  END w0_wd_in[399]
  PIN w0_wd_in[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 438.865 0.000 438.935 0.140 ;
    END
  END w0_wd_in[400]
  PIN w0_wd_in[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 441.905 0.000 441.975 0.140 ;
    END
  END w0_wd_in[401]
  PIN w0_wd_in[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 444.945 0.000 445.015 0.140 ;
    END
  END w0_wd_in[402]
  PIN w0_wd_in[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 447.985 0.000 448.055 0.140 ;
    END
  END w0_wd_in[403]
  PIN w0_wd_in[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 451.025 0.000 451.095 0.140 ;
    END
  END w0_wd_in[404]
  PIN w0_wd_in[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 454.065 0.000 454.135 0.140 ;
    END
  END w0_wd_in[405]
  PIN w0_wd_in[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 457.105 0.000 457.175 0.140 ;
    END
  END w0_wd_in[406]
  PIN w0_wd_in[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 460.145 0.000 460.215 0.140 ;
    END
  END w0_wd_in[407]
  PIN w0_wd_in[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 463.185 0.000 463.255 0.140 ;
    END
  END w0_wd_in[408]
  PIN w0_wd_in[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 466.225 0.000 466.295 0.140 ;
    END
  END w0_wd_in[409]
  PIN w0_wd_in[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 469.265 0.000 469.335 0.140 ;
    END
  END w0_wd_in[410]
  PIN w0_wd_in[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 472.305 0.000 472.375 0.140 ;
    END
  END w0_wd_in[411]
  PIN w0_wd_in[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 475.345 0.000 475.415 0.140 ;
    END
  END w0_wd_in[412]
  PIN w0_wd_in[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 478.385 0.000 478.455 0.140 ;
    END
  END w0_wd_in[413]
  PIN w0_wd_in[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 481.425 0.000 481.495 0.140 ;
    END
  END w0_wd_in[414]
  PIN w0_wd_in[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 484.465 0.000 484.535 0.140 ;
    END
  END w0_wd_in[415]
  PIN w0_wd_in[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 487.505 0.000 487.575 0.140 ;
    END
  END w0_wd_in[416]
  PIN w0_wd_in[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 490.545 0.000 490.615 0.140 ;
    END
  END w0_wd_in[417]
  PIN w0_wd_in[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 493.585 0.000 493.655 0.140 ;
    END
  END w0_wd_in[418]
  PIN w0_wd_in[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 496.625 0.000 496.695 0.140 ;
    END
  END w0_wd_in[419]
  PIN w0_wd_in[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 499.665 0.000 499.735 0.140 ;
    END
  END w0_wd_in[420]
  PIN w0_wd_in[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 502.705 0.000 502.775 0.140 ;
    END
  END w0_wd_in[421]
  PIN w0_wd_in[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 505.745 0.000 505.815 0.140 ;
    END
  END w0_wd_in[422]
  PIN w0_wd_in[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 508.785 0.000 508.855 0.140 ;
    END
  END w0_wd_in[423]
  PIN w0_wd_in[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 511.825 0.000 511.895 0.140 ;
    END
  END w0_wd_in[424]
  PIN w0_wd_in[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 514.865 0.000 514.935 0.140 ;
    END
  END w0_wd_in[425]
  PIN w0_wd_in[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 517.905 0.000 517.975 0.140 ;
    END
  END w0_wd_in[426]
  PIN w0_wd_in[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 520.945 0.000 521.015 0.140 ;
    END
  END w0_wd_in[427]
  PIN w0_wd_in[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 523.985 0.000 524.055 0.140 ;
    END
  END w0_wd_in[428]
  PIN w0_wd_in[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 527.025 0.000 527.095 0.140 ;
    END
  END w0_wd_in[429]
  PIN w0_wd_in[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 530.065 0.000 530.135 0.140 ;
    END
  END w0_wd_in[430]
  PIN w0_wd_in[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 533.105 0.000 533.175 0.140 ;
    END
  END w0_wd_in[431]
  PIN w0_wd_in[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 536.145 0.000 536.215 0.140 ;
    END
  END w0_wd_in[432]
  PIN w0_wd_in[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 539.185 0.000 539.255 0.140 ;
    END
  END w0_wd_in[433]
  PIN w0_wd_in[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 542.225 0.000 542.295 0.140 ;
    END
  END w0_wd_in[434]
  PIN w0_wd_in[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 545.265 0.000 545.335 0.140 ;
    END
  END w0_wd_in[435]
  PIN w0_wd_in[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 548.305 0.000 548.375 0.140 ;
    END
  END w0_wd_in[436]
  PIN w0_wd_in[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 551.345 0.000 551.415 0.140 ;
    END
  END w0_wd_in[437]
  PIN w0_wd_in[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 554.385 0.000 554.455 0.140 ;
    END
  END w0_wd_in[438]
  PIN w0_wd_in[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 557.425 0.000 557.495 0.140 ;
    END
  END w0_wd_in[439]
  PIN w0_wd_in[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 560.465 0.000 560.535 0.140 ;
    END
  END w0_wd_in[440]
  PIN w0_wd_in[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 563.505 0.000 563.575 0.140 ;
    END
  END w0_wd_in[441]
  PIN w0_wd_in[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 566.545 0.000 566.615 0.140 ;
    END
  END w0_wd_in[442]
  PIN w0_wd_in[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 569.585 0.000 569.655 0.140 ;
    END
  END w0_wd_in[443]
  PIN w0_wd_in[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 572.625 0.000 572.695 0.140 ;
    END
  END w0_wd_in[444]
  PIN w0_wd_in[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 575.665 0.000 575.735 0.140 ;
    END
  END w0_wd_in[445]
  PIN w0_wd_in[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 578.705 0.000 578.775 0.140 ;
    END
  END w0_wd_in[446]
  PIN w0_wd_in[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 581.745 0.000 581.815 0.140 ;
    END
  END w0_wd_in[447]
  PIN w0_wd_in[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 584.785 0.000 584.855 0.140 ;
    END
  END w0_wd_in[448]
  PIN w0_wd_in[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 587.825 0.000 587.895 0.140 ;
    END
  END w0_wd_in[449]
  PIN w0_wd_in[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 590.865 0.000 590.935 0.140 ;
    END
  END w0_wd_in[450]
  PIN w0_wd_in[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 593.905 0.000 593.975 0.140 ;
    END
  END w0_wd_in[451]
  PIN w0_wd_in[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 596.945 0.000 597.015 0.140 ;
    END
  END w0_wd_in[452]
  PIN w0_wd_in[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 599.985 0.000 600.055 0.140 ;
    END
  END w0_wd_in[453]
  PIN w0_wd_in[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 603.025 0.000 603.095 0.140 ;
    END
  END w0_wd_in[454]
  PIN w0_wd_in[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 606.065 0.000 606.135 0.140 ;
    END
  END w0_wd_in[455]
  PIN w0_wd_in[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 609.105 0.000 609.175 0.140 ;
    END
  END w0_wd_in[456]
  PIN w0_wd_in[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 612.145 0.000 612.215 0.140 ;
    END
  END w0_wd_in[457]
  PIN w0_wd_in[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 615.185 0.000 615.255 0.140 ;
    END
  END w0_wd_in[458]
  PIN w0_wd_in[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 618.225 0.000 618.295 0.140 ;
    END
  END w0_wd_in[459]
  PIN w0_wd_in[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 621.265 0.000 621.335 0.140 ;
    END
  END w0_wd_in[460]
  PIN w0_wd_in[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 624.305 0.000 624.375 0.140 ;
    END
  END w0_wd_in[461]
  PIN w0_wd_in[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 627.345 0.000 627.415 0.140 ;
    END
  END w0_wd_in[462]
  PIN w0_wd_in[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 630.385 0.000 630.455 0.140 ;
    END
  END w0_wd_in[463]
  PIN w0_wd_in[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 633.425 0.000 633.495 0.140 ;
    END
  END w0_wd_in[464]
  PIN w0_wd_in[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 636.465 0.000 636.535 0.140 ;
    END
  END w0_wd_in[465]
  PIN w0_wd_in[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 639.505 0.000 639.575 0.140 ;
    END
  END w0_wd_in[466]
  PIN w0_wd_in[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 642.545 0.000 642.615 0.140 ;
    END
  END w0_wd_in[467]
  PIN w0_wd_in[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 645.585 0.000 645.655 0.140 ;
    END
  END w0_wd_in[468]
  PIN w0_wd_in[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 648.625 0.000 648.695 0.140 ;
    END
  END w0_wd_in[469]
  PIN w0_wd_in[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 651.665 0.000 651.735 0.140 ;
    END
  END w0_wd_in[470]
  PIN w0_wd_in[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 654.705 0.000 654.775 0.140 ;
    END
  END w0_wd_in[471]
  PIN w0_wd_in[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 657.745 0.000 657.815 0.140 ;
    END
  END w0_wd_in[472]
  PIN w0_wd_in[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 660.785 0.000 660.855 0.140 ;
    END
  END w0_wd_in[473]
  PIN w0_wd_in[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 663.825 0.000 663.895 0.140 ;
    END
  END w0_wd_in[474]
  PIN w0_wd_in[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 666.865 0.000 666.935 0.140 ;
    END
  END w0_wd_in[475]
  PIN w0_wd_in[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 669.905 0.000 669.975 0.140 ;
    END
  END w0_wd_in[476]
  PIN w0_wd_in[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 672.945 0.000 673.015 0.140 ;
    END
  END w0_wd_in[477]
  PIN w0_wd_in[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 675.985 0.000 676.055 0.140 ;
    END
  END w0_wd_in[478]
  PIN w0_wd_in[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 679.025 0.000 679.095 0.140 ;
    END
  END w0_wd_in[479]
  PIN w0_wd_in[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 682.065 0.000 682.135 0.140 ;
    END
  END w0_wd_in[480]
  PIN w0_wd_in[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 685.105 0.000 685.175 0.140 ;
    END
  END w0_wd_in[481]
  PIN w0_wd_in[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 688.145 0.000 688.215 0.140 ;
    END
  END w0_wd_in[482]
  PIN w0_wd_in[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 691.185 0.000 691.255 0.140 ;
    END
  END w0_wd_in[483]
  PIN w0_wd_in[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 694.225 0.000 694.295 0.140 ;
    END
  END w0_wd_in[484]
  PIN w0_wd_in[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 697.265 0.000 697.335 0.140 ;
    END
  END w0_wd_in[485]
  PIN w0_wd_in[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 700.305 0.000 700.375 0.140 ;
    END
  END w0_wd_in[486]
  PIN w0_wd_in[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 703.345 0.000 703.415 0.140 ;
    END
  END w0_wd_in[487]
  PIN w0_wd_in[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 706.385 0.000 706.455 0.140 ;
    END
  END w0_wd_in[488]
  PIN w0_wd_in[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 709.425 0.000 709.495 0.140 ;
    END
  END w0_wd_in[489]
  PIN w0_wd_in[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 712.465 0.000 712.535 0.140 ;
    END
  END w0_wd_in[490]
  PIN w0_wd_in[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 715.505 0.000 715.575 0.140 ;
    END
  END w0_wd_in[491]
  PIN w0_wd_in[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 718.545 0.000 718.615 0.140 ;
    END
  END w0_wd_in[492]
  PIN w0_wd_in[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 721.585 0.000 721.655 0.140 ;
    END
  END w0_wd_in[493]
  PIN w0_wd_in[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 724.625 0.000 724.695 0.140 ;
    END
  END w0_wd_in[494]
  PIN w0_wd_in[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 727.665 0.000 727.735 0.140 ;
    END
  END w0_wd_in[495]
  PIN w0_wd_in[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 730.705 0.000 730.775 0.140 ;
    END
  END w0_wd_in[496]
  PIN w0_wd_in[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 733.745 0.000 733.815 0.140 ;
    END
  END w0_wd_in[497]
  PIN w0_wd_in[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 736.785 0.000 736.855 0.140 ;
    END
  END w0_wd_in[498]
  PIN w0_wd_in[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 739.825 0.000 739.895 0.140 ;
    END
  END w0_wd_in[499]
  PIN w0_wd_in[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 742.865 0.000 742.935 0.140 ;
    END
  END w0_wd_in[500]
  PIN w0_wd_in[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 745.905 0.000 745.975 0.140 ;
    END
  END w0_wd_in[501]
  PIN w0_wd_in[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 748.945 0.000 749.015 0.140 ;
    END
  END w0_wd_in[502]
  PIN w0_wd_in[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 751.985 0.000 752.055 0.140 ;
    END
  END w0_wd_in[503]
  PIN w0_wd_in[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 755.025 0.000 755.095 0.140 ;
    END
  END w0_wd_in[504]
  PIN w0_wd_in[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 758.065 0.000 758.135 0.140 ;
    END
  END w0_wd_in[505]
  PIN w0_wd_in[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 761.105 0.000 761.175 0.140 ;
    END
  END w0_wd_in[506]
  PIN w0_wd_in[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 764.145 0.000 764.215 0.140 ;
    END
  END w0_wd_in[507]
  PIN w0_wd_in[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 767.185 0.000 767.255 0.140 ;
    END
  END w0_wd_in[508]
  PIN w0_wd_in[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 770.225 0.000 770.295 0.140 ;
    END
  END w0_wd_in[509]
  PIN w0_wd_in[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 773.265 0.000 773.335 0.140 ;
    END
  END w0_wd_in[510]
  PIN w0_wd_in[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 776.305 0.000 776.375 0.140 ;
    END
  END w0_wd_in[511]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 779.345 0.000 779.415 0.140 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 782.385 0.000 782.455 0.140 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 785.425 0.000 785.495 0.140 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 788.465 0.000 788.535 0.140 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 791.505 0.000 791.575 0.140 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 794.545 0.000 794.615 0.140 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 797.585 0.000 797.655 0.140 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 800.625 0.000 800.695 0.140 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 803.665 0.000 803.735 0.140 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 806.705 0.000 806.775 0.140 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 809.745 0.000 809.815 0.140 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 812.785 0.000 812.855 0.140 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 815.825 0.000 815.895 0.140 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 818.865 0.000 818.935 0.140 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 821.905 0.000 821.975 0.140 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 824.945 0.000 825.015 0.140 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 827.985 0.000 828.055 0.140 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 831.025 0.000 831.095 0.140 ;
    END
  END r0_rd_out[17]
  PIN r0_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 834.065 0.000 834.135 0.140 ;
    END
  END r0_rd_out[18]
  PIN r0_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 837.105 0.000 837.175 0.140 ;
    END
  END r0_rd_out[19]
  PIN r0_rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 840.145 0.000 840.215 0.140 ;
    END
  END r0_rd_out[20]
  PIN r0_rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 843.185 0.000 843.255 0.140 ;
    END
  END r0_rd_out[21]
  PIN r0_rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 846.225 0.000 846.295 0.140 ;
    END
  END r0_rd_out[22]
  PIN r0_rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 849.265 0.000 849.335 0.140 ;
    END
  END r0_rd_out[23]
  PIN r0_rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 852.305 0.000 852.375 0.140 ;
    END
  END r0_rd_out[24]
  PIN r0_rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 855.345 0.000 855.415 0.140 ;
    END
  END r0_rd_out[25]
  PIN r0_rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 858.385 0.000 858.455 0.140 ;
    END
  END r0_rd_out[26]
  PIN r0_rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 861.425 0.000 861.495 0.140 ;
    END
  END r0_rd_out[27]
  PIN r0_rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 864.465 0.000 864.535 0.140 ;
    END
  END r0_rd_out[28]
  PIN r0_rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 867.505 0.000 867.575 0.140 ;
    END
  END r0_rd_out[29]
  PIN r0_rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 870.545 0.000 870.615 0.140 ;
    END
  END r0_rd_out[30]
  PIN r0_rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 873.585 0.000 873.655 0.140 ;
    END
  END r0_rd_out[31]
  PIN r0_rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 876.625 0.000 876.695 0.140 ;
    END
  END r0_rd_out[32]
  PIN r0_rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 879.665 0.000 879.735 0.140 ;
    END
  END r0_rd_out[33]
  PIN r0_rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 882.705 0.000 882.775 0.140 ;
    END
  END r0_rd_out[34]
  PIN r0_rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 885.745 0.000 885.815 0.140 ;
    END
  END r0_rd_out[35]
  PIN r0_rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 888.785 0.000 888.855 0.140 ;
    END
  END r0_rd_out[36]
  PIN r0_rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 891.825 0.000 891.895 0.140 ;
    END
  END r0_rd_out[37]
  PIN r0_rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 894.865 0.000 894.935 0.140 ;
    END
  END r0_rd_out[38]
  PIN r0_rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 897.905 0.000 897.975 0.140 ;
    END
  END r0_rd_out[39]
  PIN r0_rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 900.945 0.000 901.015 0.140 ;
    END
  END r0_rd_out[40]
  PIN r0_rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 903.985 0.000 904.055 0.140 ;
    END
  END r0_rd_out[41]
  PIN r0_rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 907.025 0.000 907.095 0.140 ;
    END
  END r0_rd_out[42]
  PIN r0_rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 910.065 0.000 910.135 0.140 ;
    END
  END r0_rd_out[43]
  PIN r0_rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 913.105 0.000 913.175 0.140 ;
    END
  END r0_rd_out[44]
  PIN r0_rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 916.145 0.000 916.215 0.140 ;
    END
  END r0_rd_out[45]
  PIN r0_rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 919.185 0.000 919.255 0.140 ;
    END
  END r0_rd_out[46]
  PIN r0_rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 922.225 0.000 922.295 0.140 ;
    END
  END r0_rd_out[47]
  PIN r0_rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 925.265 0.000 925.335 0.140 ;
    END
  END r0_rd_out[48]
  PIN r0_rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 928.305 0.000 928.375 0.140 ;
    END
  END r0_rd_out[49]
  PIN r0_rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 931.345 0.000 931.415 0.140 ;
    END
  END r0_rd_out[50]
  PIN r0_rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 934.385 0.000 934.455 0.140 ;
    END
  END r0_rd_out[51]
  PIN r0_rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 937.425 0.000 937.495 0.140 ;
    END
  END r0_rd_out[52]
  PIN r0_rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 940.465 0.000 940.535 0.140 ;
    END
  END r0_rd_out[53]
  PIN r0_rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 943.505 0.000 943.575 0.140 ;
    END
  END r0_rd_out[54]
  PIN r0_rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 946.545 0.000 946.615 0.140 ;
    END
  END r0_rd_out[55]
  PIN r0_rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 949.585 0.000 949.655 0.140 ;
    END
  END r0_rd_out[56]
  PIN r0_rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 952.625 0.000 952.695 0.140 ;
    END
  END r0_rd_out[57]
  PIN r0_rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 955.665 0.000 955.735 0.140 ;
    END
  END r0_rd_out[58]
  PIN r0_rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 958.705 0.000 958.775 0.140 ;
    END
  END r0_rd_out[59]
  PIN r0_rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 961.745 0.000 961.815 0.140 ;
    END
  END r0_rd_out[60]
  PIN r0_rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 964.785 0.000 964.855 0.140 ;
    END
  END r0_rd_out[61]
  PIN r0_rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 967.825 0.000 967.895 0.140 ;
    END
  END r0_rd_out[62]
  PIN r0_rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 970.865 0.000 970.935 0.140 ;
    END
  END r0_rd_out[63]
  PIN r0_rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 973.905 0.000 973.975 0.140 ;
    END
  END r0_rd_out[64]
  PIN r0_rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 976.945 0.000 977.015 0.140 ;
    END
  END r0_rd_out[65]
  PIN r0_rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 979.985 0.000 980.055 0.140 ;
    END
  END r0_rd_out[66]
  PIN r0_rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 983.025 0.000 983.095 0.140 ;
    END
  END r0_rd_out[67]
  PIN r0_rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 986.065 0.000 986.135 0.140 ;
    END
  END r0_rd_out[68]
  PIN r0_rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 989.105 0.000 989.175 0.140 ;
    END
  END r0_rd_out[69]
  PIN r0_rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 992.145 0.000 992.215 0.140 ;
    END
  END r0_rd_out[70]
  PIN r0_rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 995.185 0.000 995.255 0.140 ;
    END
  END r0_rd_out[71]
  PIN r0_rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 998.225 0.000 998.295 0.140 ;
    END
  END r0_rd_out[72]
  PIN r0_rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1001.265 0.000 1001.335 0.140 ;
    END
  END r0_rd_out[73]
  PIN r0_rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1004.305 0.000 1004.375 0.140 ;
    END
  END r0_rd_out[74]
  PIN r0_rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1007.345 0.000 1007.415 0.140 ;
    END
  END r0_rd_out[75]
  PIN r0_rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1010.385 0.000 1010.455 0.140 ;
    END
  END r0_rd_out[76]
  PIN r0_rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1013.425 0.000 1013.495 0.140 ;
    END
  END r0_rd_out[77]
  PIN r0_rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1016.465 0.000 1016.535 0.140 ;
    END
  END r0_rd_out[78]
  PIN r0_rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1019.505 0.000 1019.575 0.140 ;
    END
  END r0_rd_out[79]
  PIN r0_rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1022.545 0.000 1022.615 0.140 ;
    END
  END r0_rd_out[80]
  PIN r0_rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1025.585 0.000 1025.655 0.140 ;
    END
  END r0_rd_out[81]
  PIN r0_rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1028.625 0.000 1028.695 0.140 ;
    END
  END r0_rd_out[82]
  PIN r0_rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1031.665 0.000 1031.735 0.140 ;
    END
  END r0_rd_out[83]
  PIN r0_rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1034.705 0.000 1034.775 0.140 ;
    END
  END r0_rd_out[84]
  PIN r0_rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1037.745 0.000 1037.815 0.140 ;
    END
  END r0_rd_out[85]
  PIN r0_rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1040.785 0.000 1040.855 0.140 ;
    END
  END r0_rd_out[86]
  PIN r0_rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1043.825 0.000 1043.895 0.140 ;
    END
  END r0_rd_out[87]
  PIN r0_rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1046.865 0.000 1046.935 0.140 ;
    END
  END r0_rd_out[88]
  PIN r0_rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1049.905 0.000 1049.975 0.140 ;
    END
  END r0_rd_out[89]
  PIN r0_rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1052.945 0.000 1053.015 0.140 ;
    END
  END r0_rd_out[90]
  PIN r0_rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1055.985 0.000 1056.055 0.140 ;
    END
  END r0_rd_out[91]
  PIN r0_rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1059.025 0.000 1059.095 0.140 ;
    END
  END r0_rd_out[92]
  PIN r0_rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1062.065 0.000 1062.135 0.140 ;
    END
  END r0_rd_out[93]
  PIN r0_rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1065.105 0.000 1065.175 0.140 ;
    END
  END r0_rd_out[94]
  PIN r0_rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1068.145 0.000 1068.215 0.140 ;
    END
  END r0_rd_out[95]
  PIN r0_rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1071.185 0.000 1071.255 0.140 ;
    END
  END r0_rd_out[96]
  PIN r0_rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1074.225 0.000 1074.295 0.140 ;
    END
  END r0_rd_out[97]
  PIN r0_rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1077.265 0.000 1077.335 0.140 ;
    END
  END r0_rd_out[98]
  PIN r0_rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1080.305 0.000 1080.375 0.140 ;
    END
  END r0_rd_out[99]
  PIN r0_rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1083.345 0.000 1083.415 0.140 ;
    END
  END r0_rd_out[100]
  PIN r0_rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1086.385 0.000 1086.455 0.140 ;
    END
  END r0_rd_out[101]
  PIN r0_rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1089.425 0.000 1089.495 0.140 ;
    END
  END r0_rd_out[102]
  PIN r0_rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1092.465 0.000 1092.535 0.140 ;
    END
  END r0_rd_out[103]
  PIN r0_rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1095.505 0.000 1095.575 0.140 ;
    END
  END r0_rd_out[104]
  PIN r0_rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1098.545 0.000 1098.615 0.140 ;
    END
  END r0_rd_out[105]
  PIN r0_rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1101.585 0.000 1101.655 0.140 ;
    END
  END r0_rd_out[106]
  PIN r0_rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1104.625 0.000 1104.695 0.140 ;
    END
  END r0_rd_out[107]
  PIN r0_rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1107.665 0.000 1107.735 0.140 ;
    END
  END r0_rd_out[108]
  PIN r0_rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1110.705 0.000 1110.775 0.140 ;
    END
  END r0_rd_out[109]
  PIN r0_rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1113.745 0.000 1113.815 0.140 ;
    END
  END r0_rd_out[110]
  PIN r0_rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1116.785 0.000 1116.855 0.140 ;
    END
  END r0_rd_out[111]
  PIN r0_rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1119.825 0.000 1119.895 0.140 ;
    END
  END r0_rd_out[112]
  PIN r0_rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1122.865 0.000 1122.935 0.140 ;
    END
  END r0_rd_out[113]
  PIN r0_rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1125.905 0.000 1125.975 0.140 ;
    END
  END r0_rd_out[114]
  PIN r0_rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1128.945 0.000 1129.015 0.140 ;
    END
  END r0_rd_out[115]
  PIN r0_rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1131.985 0.000 1132.055 0.140 ;
    END
  END r0_rd_out[116]
  PIN r0_rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1135.025 0.000 1135.095 0.140 ;
    END
  END r0_rd_out[117]
  PIN r0_rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1138.065 0.000 1138.135 0.140 ;
    END
  END r0_rd_out[118]
  PIN r0_rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1141.105 0.000 1141.175 0.140 ;
    END
  END r0_rd_out[119]
  PIN r0_rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1144.145 0.000 1144.215 0.140 ;
    END
  END r0_rd_out[120]
  PIN r0_rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1147.185 0.000 1147.255 0.140 ;
    END
  END r0_rd_out[121]
  PIN r0_rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1150.225 0.000 1150.295 0.140 ;
    END
  END r0_rd_out[122]
  PIN r0_rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1153.265 0.000 1153.335 0.140 ;
    END
  END r0_rd_out[123]
  PIN r0_rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1156.305 0.000 1156.375 0.140 ;
    END
  END r0_rd_out[124]
  PIN r0_rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1159.345 0.000 1159.415 0.140 ;
    END
  END r0_rd_out[125]
  PIN r0_rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1162.385 0.000 1162.455 0.140 ;
    END
  END r0_rd_out[126]
  PIN r0_rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1165.425 0.000 1165.495 0.140 ;
    END
  END r0_rd_out[127]
  PIN r0_rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1168.465 0.000 1168.535 0.140 ;
    END
  END r0_rd_out[128]
  PIN r0_rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1171.505 0.000 1171.575 0.140 ;
    END
  END r0_rd_out[129]
  PIN r0_rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1174.545 0.000 1174.615 0.140 ;
    END
  END r0_rd_out[130]
  PIN r0_rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1177.585 0.000 1177.655 0.140 ;
    END
  END r0_rd_out[131]
  PIN r0_rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1180.625 0.000 1180.695 0.140 ;
    END
  END r0_rd_out[132]
  PIN r0_rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1183.665 0.000 1183.735 0.140 ;
    END
  END r0_rd_out[133]
  PIN r0_rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1186.705 0.000 1186.775 0.140 ;
    END
  END r0_rd_out[134]
  PIN r0_rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1189.745 0.000 1189.815 0.140 ;
    END
  END r0_rd_out[135]
  PIN r0_rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1192.785 0.000 1192.855 0.140 ;
    END
  END r0_rd_out[136]
  PIN r0_rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1195.825 0.000 1195.895 0.140 ;
    END
  END r0_rd_out[137]
  PIN r0_rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1198.865 0.000 1198.935 0.140 ;
    END
  END r0_rd_out[138]
  PIN r0_rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1201.905 0.000 1201.975 0.140 ;
    END
  END r0_rd_out[139]
  PIN r0_rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1204.945 0.000 1205.015 0.140 ;
    END
  END r0_rd_out[140]
  PIN r0_rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1207.985 0.000 1208.055 0.140 ;
    END
  END r0_rd_out[141]
  PIN r0_rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1211.025 0.000 1211.095 0.140 ;
    END
  END r0_rd_out[142]
  PIN r0_rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1214.065 0.000 1214.135 0.140 ;
    END
  END r0_rd_out[143]
  PIN r0_rd_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1217.105 0.000 1217.175 0.140 ;
    END
  END r0_rd_out[144]
  PIN r0_rd_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1220.145 0.000 1220.215 0.140 ;
    END
  END r0_rd_out[145]
  PIN r0_rd_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1223.185 0.000 1223.255 0.140 ;
    END
  END r0_rd_out[146]
  PIN r0_rd_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1226.225 0.000 1226.295 0.140 ;
    END
  END r0_rd_out[147]
  PIN r0_rd_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1229.265 0.000 1229.335 0.140 ;
    END
  END r0_rd_out[148]
  PIN r0_rd_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1232.305 0.000 1232.375 0.140 ;
    END
  END r0_rd_out[149]
  PIN r0_rd_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1235.345 0.000 1235.415 0.140 ;
    END
  END r0_rd_out[150]
  PIN r0_rd_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1238.385 0.000 1238.455 0.140 ;
    END
  END r0_rd_out[151]
  PIN r0_rd_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1241.425 0.000 1241.495 0.140 ;
    END
  END r0_rd_out[152]
  PIN r0_rd_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1244.465 0.000 1244.535 0.140 ;
    END
  END r0_rd_out[153]
  PIN r0_rd_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1247.505 0.000 1247.575 0.140 ;
    END
  END r0_rd_out[154]
  PIN r0_rd_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1250.545 0.000 1250.615 0.140 ;
    END
  END r0_rd_out[155]
  PIN r0_rd_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1253.585 0.000 1253.655 0.140 ;
    END
  END r0_rd_out[156]
  PIN r0_rd_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1256.625 0.000 1256.695 0.140 ;
    END
  END r0_rd_out[157]
  PIN r0_rd_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1259.665 0.000 1259.735 0.140 ;
    END
  END r0_rd_out[158]
  PIN r0_rd_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1262.705 0.000 1262.775 0.140 ;
    END
  END r0_rd_out[159]
  PIN r0_rd_out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1265.745 0.000 1265.815 0.140 ;
    END
  END r0_rd_out[160]
  PIN r0_rd_out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1268.785 0.000 1268.855 0.140 ;
    END
  END r0_rd_out[161]
  PIN r0_rd_out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1271.825 0.000 1271.895 0.140 ;
    END
  END r0_rd_out[162]
  PIN r0_rd_out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1274.865 0.000 1274.935 0.140 ;
    END
  END r0_rd_out[163]
  PIN r0_rd_out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1277.905 0.000 1277.975 0.140 ;
    END
  END r0_rd_out[164]
  PIN r0_rd_out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1280.945 0.000 1281.015 0.140 ;
    END
  END r0_rd_out[165]
  PIN r0_rd_out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1283.985 0.000 1284.055 0.140 ;
    END
  END r0_rd_out[166]
  PIN r0_rd_out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1287.025 0.000 1287.095 0.140 ;
    END
  END r0_rd_out[167]
  PIN r0_rd_out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1290.065 0.000 1290.135 0.140 ;
    END
  END r0_rd_out[168]
  PIN r0_rd_out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1293.105 0.000 1293.175 0.140 ;
    END
  END r0_rd_out[169]
  PIN r0_rd_out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1296.145 0.000 1296.215 0.140 ;
    END
  END r0_rd_out[170]
  PIN r0_rd_out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1299.185 0.000 1299.255 0.140 ;
    END
  END r0_rd_out[171]
  PIN r0_rd_out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1302.225 0.000 1302.295 0.140 ;
    END
  END r0_rd_out[172]
  PIN r0_rd_out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1305.265 0.000 1305.335 0.140 ;
    END
  END r0_rd_out[173]
  PIN r0_rd_out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1308.305 0.000 1308.375 0.140 ;
    END
  END r0_rd_out[174]
  PIN r0_rd_out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1311.345 0.000 1311.415 0.140 ;
    END
  END r0_rd_out[175]
  PIN r0_rd_out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1314.385 0.000 1314.455 0.140 ;
    END
  END r0_rd_out[176]
  PIN r0_rd_out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1317.425 0.000 1317.495 0.140 ;
    END
  END r0_rd_out[177]
  PIN r0_rd_out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1320.465 0.000 1320.535 0.140 ;
    END
  END r0_rd_out[178]
  PIN r0_rd_out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1323.505 0.000 1323.575 0.140 ;
    END
  END r0_rd_out[179]
  PIN r0_rd_out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1326.545 0.000 1326.615 0.140 ;
    END
  END r0_rd_out[180]
  PIN r0_rd_out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1329.585 0.000 1329.655 0.140 ;
    END
  END r0_rd_out[181]
  PIN r0_rd_out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1332.625 0.000 1332.695 0.140 ;
    END
  END r0_rd_out[182]
  PIN r0_rd_out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1335.665 0.000 1335.735 0.140 ;
    END
  END r0_rd_out[183]
  PIN r0_rd_out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1338.705 0.000 1338.775 0.140 ;
    END
  END r0_rd_out[184]
  PIN r0_rd_out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1341.745 0.000 1341.815 0.140 ;
    END
  END r0_rd_out[185]
  PIN r0_rd_out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1344.785 0.000 1344.855 0.140 ;
    END
  END r0_rd_out[186]
  PIN r0_rd_out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1347.825 0.000 1347.895 0.140 ;
    END
  END r0_rd_out[187]
  PIN r0_rd_out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1350.865 0.000 1350.935 0.140 ;
    END
  END r0_rd_out[188]
  PIN r0_rd_out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1353.905 0.000 1353.975 0.140 ;
    END
  END r0_rd_out[189]
  PIN r0_rd_out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1356.945 0.000 1357.015 0.140 ;
    END
  END r0_rd_out[190]
  PIN r0_rd_out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1359.985 0.000 1360.055 0.140 ;
    END
  END r0_rd_out[191]
  PIN r0_rd_out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1363.025 0.000 1363.095 0.140 ;
    END
  END r0_rd_out[192]
  PIN r0_rd_out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1366.065 0.000 1366.135 0.140 ;
    END
  END r0_rd_out[193]
  PIN r0_rd_out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1369.105 0.000 1369.175 0.140 ;
    END
  END r0_rd_out[194]
  PIN r0_rd_out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1372.145 0.000 1372.215 0.140 ;
    END
  END r0_rd_out[195]
  PIN r0_rd_out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1375.185 0.000 1375.255 0.140 ;
    END
  END r0_rd_out[196]
  PIN r0_rd_out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1378.225 0.000 1378.295 0.140 ;
    END
  END r0_rd_out[197]
  PIN r0_rd_out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1381.265 0.000 1381.335 0.140 ;
    END
  END r0_rd_out[198]
  PIN r0_rd_out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1384.305 0.000 1384.375 0.140 ;
    END
  END r0_rd_out[199]
  PIN r0_rd_out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1387.345 0.000 1387.415 0.140 ;
    END
  END r0_rd_out[200]
  PIN r0_rd_out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1390.385 0.000 1390.455 0.140 ;
    END
  END r0_rd_out[201]
  PIN r0_rd_out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1393.425 0.000 1393.495 0.140 ;
    END
  END r0_rd_out[202]
  PIN r0_rd_out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1396.465 0.000 1396.535 0.140 ;
    END
  END r0_rd_out[203]
  PIN r0_rd_out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1399.505 0.000 1399.575 0.140 ;
    END
  END r0_rd_out[204]
  PIN r0_rd_out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1402.545 0.000 1402.615 0.140 ;
    END
  END r0_rd_out[205]
  PIN r0_rd_out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1405.585 0.000 1405.655 0.140 ;
    END
  END r0_rd_out[206]
  PIN r0_rd_out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1408.625 0.000 1408.695 0.140 ;
    END
  END r0_rd_out[207]
  PIN r0_rd_out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1411.665 0.000 1411.735 0.140 ;
    END
  END r0_rd_out[208]
  PIN r0_rd_out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1414.705 0.000 1414.775 0.140 ;
    END
  END r0_rd_out[209]
  PIN r0_rd_out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1417.745 0.000 1417.815 0.140 ;
    END
  END r0_rd_out[210]
  PIN r0_rd_out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1420.785 0.000 1420.855 0.140 ;
    END
  END r0_rd_out[211]
  PIN r0_rd_out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1423.825 0.000 1423.895 0.140 ;
    END
  END r0_rd_out[212]
  PIN r0_rd_out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1426.865 0.000 1426.935 0.140 ;
    END
  END r0_rd_out[213]
  PIN r0_rd_out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1429.905 0.000 1429.975 0.140 ;
    END
  END r0_rd_out[214]
  PIN r0_rd_out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1432.945 0.000 1433.015 0.140 ;
    END
  END r0_rd_out[215]
  PIN r0_rd_out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1435.985 0.000 1436.055 0.140 ;
    END
  END r0_rd_out[216]
  PIN r0_rd_out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1439.025 0.000 1439.095 0.140 ;
    END
  END r0_rd_out[217]
  PIN r0_rd_out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1442.065 0.000 1442.135 0.140 ;
    END
  END r0_rd_out[218]
  PIN r0_rd_out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1445.105 0.000 1445.175 0.140 ;
    END
  END r0_rd_out[219]
  PIN r0_rd_out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1448.145 0.000 1448.215 0.140 ;
    END
  END r0_rd_out[220]
  PIN r0_rd_out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1451.185 0.000 1451.255 0.140 ;
    END
  END r0_rd_out[221]
  PIN r0_rd_out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1454.225 0.000 1454.295 0.140 ;
    END
  END r0_rd_out[222]
  PIN r0_rd_out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1457.265 0.000 1457.335 0.140 ;
    END
  END r0_rd_out[223]
  PIN r0_rd_out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1460.305 0.000 1460.375 0.140 ;
    END
  END r0_rd_out[224]
  PIN r0_rd_out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1463.345 0.000 1463.415 0.140 ;
    END
  END r0_rd_out[225]
  PIN r0_rd_out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1466.385 0.000 1466.455 0.140 ;
    END
  END r0_rd_out[226]
  PIN r0_rd_out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1469.425 0.000 1469.495 0.140 ;
    END
  END r0_rd_out[227]
  PIN r0_rd_out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1472.465 0.000 1472.535 0.140 ;
    END
  END r0_rd_out[228]
  PIN r0_rd_out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1475.505 0.000 1475.575 0.140 ;
    END
  END r0_rd_out[229]
  PIN r0_rd_out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1478.545 0.000 1478.615 0.140 ;
    END
  END r0_rd_out[230]
  PIN r0_rd_out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1481.585 0.000 1481.655 0.140 ;
    END
  END r0_rd_out[231]
  PIN r0_rd_out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1484.625 0.000 1484.695 0.140 ;
    END
  END r0_rd_out[232]
  PIN r0_rd_out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1487.665 0.000 1487.735 0.140 ;
    END
  END r0_rd_out[233]
  PIN r0_rd_out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1490.705 0.000 1490.775 0.140 ;
    END
  END r0_rd_out[234]
  PIN r0_rd_out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1493.745 0.000 1493.815 0.140 ;
    END
  END r0_rd_out[235]
  PIN r0_rd_out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1496.785 0.000 1496.855 0.140 ;
    END
  END r0_rd_out[236]
  PIN r0_rd_out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1499.825 0.000 1499.895 0.140 ;
    END
  END r0_rd_out[237]
  PIN r0_rd_out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1502.865 0.000 1502.935 0.140 ;
    END
  END r0_rd_out[238]
  PIN r0_rd_out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1505.905 0.000 1505.975 0.140 ;
    END
  END r0_rd_out[239]
  PIN r0_rd_out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1508.945 0.000 1509.015 0.140 ;
    END
  END r0_rd_out[240]
  PIN r0_rd_out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1511.985 0.000 1512.055 0.140 ;
    END
  END r0_rd_out[241]
  PIN r0_rd_out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1515.025 0.000 1515.095 0.140 ;
    END
  END r0_rd_out[242]
  PIN r0_rd_out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1518.065 0.000 1518.135 0.140 ;
    END
  END r0_rd_out[243]
  PIN r0_rd_out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1521.105 0.000 1521.175 0.140 ;
    END
  END r0_rd_out[244]
  PIN r0_rd_out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1524.145 0.000 1524.215 0.140 ;
    END
  END r0_rd_out[245]
  PIN r0_rd_out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1527.185 0.000 1527.255 0.140 ;
    END
  END r0_rd_out[246]
  PIN r0_rd_out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1530.225 0.000 1530.295 0.140 ;
    END
  END r0_rd_out[247]
  PIN r0_rd_out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1533.265 0.000 1533.335 0.140 ;
    END
  END r0_rd_out[248]
  PIN r0_rd_out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1536.305 0.000 1536.375 0.140 ;
    END
  END r0_rd_out[249]
  PIN r0_rd_out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1539.345 0.000 1539.415 0.140 ;
    END
  END r0_rd_out[250]
  PIN r0_rd_out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1542.385 0.000 1542.455 0.140 ;
    END
  END r0_rd_out[251]
  PIN r0_rd_out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1545.425 0.000 1545.495 0.140 ;
    END
  END r0_rd_out[252]
  PIN r0_rd_out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1548.465 0.000 1548.535 0.140 ;
    END
  END r0_rd_out[253]
  PIN r0_rd_out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1551.505 0.000 1551.575 0.140 ;
    END
  END r0_rd_out[254]
  PIN r0_rd_out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1554.545 0.000 1554.615 0.140 ;
    END
  END r0_rd_out[255]
  PIN r0_rd_out[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1.105 1511.860 1.175 1512.000 ;
    END
  END r0_rd_out[256]
  PIN r0_rd_out[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 7.185 1511.860 7.255 1512.000 ;
    END
  END r0_rd_out[257]
  PIN r0_rd_out[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 13.265 1511.860 13.335 1512.000 ;
    END
  END r0_rd_out[258]
  PIN r0_rd_out[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 19.345 1511.860 19.415 1512.000 ;
    END
  END r0_rd_out[259]
  PIN r0_rd_out[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 25.425 1511.860 25.495 1512.000 ;
    END
  END r0_rd_out[260]
  PIN r0_rd_out[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 31.505 1511.860 31.575 1512.000 ;
    END
  END r0_rd_out[261]
  PIN r0_rd_out[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 37.585 1511.860 37.655 1512.000 ;
    END
  END r0_rd_out[262]
  PIN r0_rd_out[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 43.665 1511.860 43.735 1512.000 ;
    END
  END r0_rd_out[263]
  PIN r0_rd_out[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 49.745 1511.860 49.815 1512.000 ;
    END
  END r0_rd_out[264]
  PIN r0_rd_out[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 55.825 1511.860 55.895 1512.000 ;
    END
  END r0_rd_out[265]
  PIN r0_rd_out[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 61.905 1511.860 61.975 1512.000 ;
    END
  END r0_rd_out[266]
  PIN r0_rd_out[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 67.985 1511.860 68.055 1512.000 ;
    END
  END r0_rd_out[267]
  PIN r0_rd_out[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 74.065 1511.860 74.135 1512.000 ;
    END
  END r0_rd_out[268]
  PIN r0_rd_out[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 80.145 1511.860 80.215 1512.000 ;
    END
  END r0_rd_out[269]
  PIN r0_rd_out[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 86.225 1511.860 86.295 1512.000 ;
    END
  END r0_rd_out[270]
  PIN r0_rd_out[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 92.305 1511.860 92.375 1512.000 ;
    END
  END r0_rd_out[271]
  PIN r0_rd_out[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 98.385 1511.860 98.455 1512.000 ;
    END
  END r0_rd_out[272]
  PIN r0_rd_out[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 104.465 1511.860 104.535 1512.000 ;
    END
  END r0_rd_out[273]
  PIN r0_rd_out[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 110.545 1511.860 110.615 1512.000 ;
    END
  END r0_rd_out[274]
  PIN r0_rd_out[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 116.625 1511.860 116.695 1512.000 ;
    END
  END r0_rd_out[275]
  PIN r0_rd_out[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 122.705 1511.860 122.775 1512.000 ;
    END
  END r0_rd_out[276]
  PIN r0_rd_out[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 128.785 1511.860 128.855 1512.000 ;
    END
  END r0_rd_out[277]
  PIN r0_rd_out[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 134.865 1511.860 134.935 1512.000 ;
    END
  END r0_rd_out[278]
  PIN r0_rd_out[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 140.945 1511.860 141.015 1512.000 ;
    END
  END r0_rd_out[279]
  PIN r0_rd_out[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 147.025 1511.860 147.095 1512.000 ;
    END
  END r0_rd_out[280]
  PIN r0_rd_out[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 153.105 1511.860 153.175 1512.000 ;
    END
  END r0_rd_out[281]
  PIN r0_rd_out[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 159.185 1511.860 159.255 1512.000 ;
    END
  END r0_rd_out[282]
  PIN r0_rd_out[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 165.265 1511.860 165.335 1512.000 ;
    END
  END r0_rd_out[283]
  PIN r0_rd_out[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 171.345 1511.860 171.415 1512.000 ;
    END
  END r0_rd_out[284]
  PIN r0_rd_out[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 177.425 1511.860 177.495 1512.000 ;
    END
  END r0_rd_out[285]
  PIN r0_rd_out[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 183.505 1511.860 183.575 1512.000 ;
    END
  END r0_rd_out[286]
  PIN r0_rd_out[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 189.585 1511.860 189.655 1512.000 ;
    END
  END r0_rd_out[287]
  PIN r0_rd_out[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 195.665 1511.860 195.735 1512.000 ;
    END
  END r0_rd_out[288]
  PIN r0_rd_out[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 201.745 1511.860 201.815 1512.000 ;
    END
  END r0_rd_out[289]
  PIN r0_rd_out[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 207.825 1511.860 207.895 1512.000 ;
    END
  END r0_rd_out[290]
  PIN r0_rd_out[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 213.905 1511.860 213.975 1512.000 ;
    END
  END r0_rd_out[291]
  PIN r0_rd_out[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 219.985 1511.860 220.055 1512.000 ;
    END
  END r0_rd_out[292]
  PIN r0_rd_out[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 226.065 1511.860 226.135 1512.000 ;
    END
  END r0_rd_out[293]
  PIN r0_rd_out[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 232.145 1511.860 232.215 1512.000 ;
    END
  END r0_rd_out[294]
  PIN r0_rd_out[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 238.225 1511.860 238.295 1512.000 ;
    END
  END r0_rd_out[295]
  PIN r0_rd_out[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 244.305 1511.860 244.375 1512.000 ;
    END
  END r0_rd_out[296]
  PIN r0_rd_out[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 250.385 1511.860 250.455 1512.000 ;
    END
  END r0_rd_out[297]
  PIN r0_rd_out[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 256.465 1511.860 256.535 1512.000 ;
    END
  END r0_rd_out[298]
  PIN r0_rd_out[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 262.545 1511.860 262.615 1512.000 ;
    END
  END r0_rd_out[299]
  PIN r0_rd_out[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 268.625 1511.860 268.695 1512.000 ;
    END
  END r0_rd_out[300]
  PIN r0_rd_out[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 274.705 1511.860 274.775 1512.000 ;
    END
  END r0_rd_out[301]
  PIN r0_rd_out[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 280.785 1511.860 280.855 1512.000 ;
    END
  END r0_rd_out[302]
  PIN r0_rd_out[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 286.865 1511.860 286.935 1512.000 ;
    END
  END r0_rd_out[303]
  PIN r0_rd_out[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 292.945 1511.860 293.015 1512.000 ;
    END
  END r0_rd_out[304]
  PIN r0_rd_out[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 299.025 1511.860 299.095 1512.000 ;
    END
  END r0_rd_out[305]
  PIN r0_rd_out[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 305.105 1511.860 305.175 1512.000 ;
    END
  END r0_rd_out[306]
  PIN r0_rd_out[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 311.185 1511.860 311.255 1512.000 ;
    END
  END r0_rd_out[307]
  PIN r0_rd_out[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 317.265 1511.860 317.335 1512.000 ;
    END
  END r0_rd_out[308]
  PIN r0_rd_out[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 323.345 1511.860 323.415 1512.000 ;
    END
  END r0_rd_out[309]
  PIN r0_rd_out[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 329.425 1511.860 329.495 1512.000 ;
    END
  END r0_rd_out[310]
  PIN r0_rd_out[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 335.505 1511.860 335.575 1512.000 ;
    END
  END r0_rd_out[311]
  PIN r0_rd_out[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 341.585 1511.860 341.655 1512.000 ;
    END
  END r0_rd_out[312]
  PIN r0_rd_out[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 347.665 1511.860 347.735 1512.000 ;
    END
  END r0_rd_out[313]
  PIN r0_rd_out[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 353.745 1511.860 353.815 1512.000 ;
    END
  END r0_rd_out[314]
  PIN r0_rd_out[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 359.825 1511.860 359.895 1512.000 ;
    END
  END r0_rd_out[315]
  PIN r0_rd_out[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 365.905 1511.860 365.975 1512.000 ;
    END
  END r0_rd_out[316]
  PIN r0_rd_out[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 371.985 1511.860 372.055 1512.000 ;
    END
  END r0_rd_out[317]
  PIN r0_rd_out[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 378.065 1511.860 378.135 1512.000 ;
    END
  END r0_rd_out[318]
  PIN r0_rd_out[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 384.145 1511.860 384.215 1512.000 ;
    END
  END r0_rd_out[319]
  PIN r0_rd_out[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 390.225 1511.860 390.295 1512.000 ;
    END
  END r0_rd_out[320]
  PIN r0_rd_out[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 396.305 1511.860 396.375 1512.000 ;
    END
  END r0_rd_out[321]
  PIN r0_rd_out[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 402.385 1511.860 402.455 1512.000 ;
    END
  END r0_rd_out[322]
  PIN r0_rd_out[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 408.465 1511.860 408.535 1512.000 ;
    END
  END r0_rd_out[323]
  PIN r0_rd_out[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 414.545 1511.860 414.615 1512.000 ;
    END
  END r0_rd_out[324]
  PIN r0_rd_out[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 420.625 1511.860 420.695 1512.000 ;
    END
  END r0_rd_out[325]
  PIN r0_rd_out[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 426.705 1511.860 426.775 1512.000 ;
    END
  END r0_rd_out[326]
  PIN r0_rd_out[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 432.785 1511.860 432.855 1512.000 ;
    END
  END r0_rd_out[327]
  PIN r0_rd_out[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 438.865 1511.860 438.935 1512.000 ;
    END
  END r0_rd_out[328]
  PIN r0_rd_out[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 444.945 1511.860 445.015 1512.000 ;
    END
  END r0_rd_out[329]
  PIN r0_rd_out[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 451.025 1511.860 451.095 1512.000 ;
    END
  END r0_rd_out[330]
  PIN r0_rd_out[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 457.105 1511.860 457.175 1512.000 ;
    END
  END r0_rd_out[331]
  PIN r0_rd_out[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 463.185 1511.860 463.255 1512.000 ;
    END
  END r0_rd_out[332]
  PIN r0_rd_out[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 469.265 1511.860 469.335 1512.000 ;
    END
  END r0_rd_out[333]
  PIN r0_rd_out[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 475.345 1511.860 475.415 1512.000 ;
    END
  END r0_rd_out[334]
  PIN r0_rd_out[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 481.425 1511.860 481.495 1512.000 ;
    END
  END r0_rd_out[335]
  PIN r0_rd_out[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 487.505 1511.860 487.575 1512.000 ;
    END
  END r0_rd_out[336]
  PIN r0_rd_out[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 493.585 1511.860 493.655 1512.000 ;
    END
  END r0_rd_out[337]
  PIN r0_rd_out[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 499.665 1511.860 499.735 1512.000 ;
    END
  END r0_rd_out[338]
  PIN r0_rd_out[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 505.745 1511.860 505.815 1512.000 ;
    END
  END r0_rd_out[339]
  PIN r0_rd_out[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 511.825 1511.860 511.895 1512.000 ;
    END
  END r0_rd_out[340]
  PIN r0_rd_out[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 517.905 1511.860 517.975 1512.000 ;
    END
  END r0_rd_out[341]
  PIN r0_rd_out[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 523.985 1511.860 524.055 1512.000 ;
    END
  END r0_rd_out[342]
  PIN r0_rd_out[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 530.065 1511.860 530.135 1512.000 ;
    END
  END r0_rd_out[343]
  PIN r0_rd_out[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 536.145 1511.860 536.215 1512.000 ;
    END
  END r0_rd_out[344]
  PIN r0_rd_out[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 542.225 1511.860 542.295 1512.000 ;
    END
  END r0_rd_out[345]
  PIN r0_rd_out[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 548.305 1511.860 548.375 1512.000 ;
    END
  END r0_rd_out[346]
  PIN r0_rd_out[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 554.385 1511.860 554.455 1512.000 ;
    END
  END r0_rd_out[347]
  PIN r0_rd_out[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 560.465 1511.860 560.535 1512.000 ;
    END
  END r0_rd_out[348]
  PIN r0_rd_out[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 566.545 1511.860 566.615 1512.000 ;
    END
  END r0_rd_out[349]
  PIN r0_rd_out[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 572.625 1511.860 572.695 1512.000 ;
    END
  END r0_rd_out[350]
  PIN r0_rd_out[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 578.705 1511.860 578.775 1512.000 ;
    END
  END r0_rd_out[351]
  PIN r0_rd_out[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 584.785 1511.860 584.855 1512.000 ;
    END
  END r0_rd_out[352]
  PIN r0_rd_out[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 590.865 1511.860 590.935 1512.000 ;
    END
  END r0_rd_out[353]
  PIN r0_rd_out[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 596.945 1511.860 597.015 1512.000 ;
    END
  END r0_rd_out[354]
  PIN r0_rd_out[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 603.025 1511.860 603.095 1512.000 ;
    END
  END r0_rd_out[355]
  PIN r0_rd_out[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 609.105 1511.860 609.175 1512.000 ;
    END
  END r0_rd_out[356]
  PIN r0_rd_out[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 615.185 1511.860 615.255 1512.000 ;
    END
  END r0_rd_out[357]
  PIN r0_rd_out[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 621.265 1511.860 621.335 1512.000 ;
    END
  END r0_rd_out[358]
  PIN r0_rd_out[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 627.345 1511.860 627.415 1512.000 ;
    END
  END r0_rd_out[359]
  PIN r0_rd_out[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 633.425 1511.860 633.495 1512.000 ;
    END
  END r0_rd_out[360]
  PIN r0_rd_out[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 639.505 1511.860 639.575 1512.000 ;
    END
  END r0_rd_out[361]
  PIN r0_rd_out[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 645.585 1511.860 645.655 1512.000 ;
    END
  END r0_rd_out[362]
  PIN r0_rd_out[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 651.665 1511.860 651.735 1512.000 ;
    END
  END r0_rd_out[363]
  PIN r0_rd_out[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 657.745 1511.860 657.815 1512.000 ;
    END
  END r0_rd_out[364]
  PIN r0_rd_out[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 663.825 1511.860 663.895 1512.000 ;
    END
  END r0_rd_out[365]
  PIN r0_rd_out[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 669.905 1511.860 669.975 1512.000 ;
    END
  END r0_rd_out[366]
  PIN r0_rd_out[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 675.985 1511.860 676.055 1512.000 ;
    END
  END r0_rd_out[367]
  PIN r0_rd_out[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 682.065 1511.860 682.135 1512.000 ;
    END
  END r0_rd_out[368]
  PIN r0_rd_out[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 688.145 1511.860 688.215 1512.000 ;
    END
  END r0_rd_out[369]
  PIN r0_rd_out[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 694.225 1511.860 694.295 1512.000 ;
    END
  END r0_rd_out[370]
  PIN r0_rd_out[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 700.305 1511.860 700.375 1512.000 ;
    END
  END r0_rd_out[371]
  PIN r0_rd_out[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 706.385 1511.860 706.455 1512.000 ;
    END
  END r0_rd_out[372]
  PIN r0_rd_out[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 712.465 1511.860 712.535 1512.000 ;
    END
  END r0_rd_out[373]
  PIN r0_rd_out[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 718.545 1511.860 718.615 1512.000 ;
    END
  END r0_rd_out[374]
  PIN r0_rd_out[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 724.625 1511.860 724.695 1512.000 ;
    END
  END r0_rd_out[375]
  PIN r0_rd_out[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 730.705 1511.860 730.775 1512.000 ;
    END
  END r0_rd_out[376]
  PIN r0_rd_out[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 736.785 1511.860 736.855 1512.000 ;
    END
  END r0_rd_out[377]
  PIN r0_rd_out[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 742.865 1511.860 742.935 1512.000 ;
    END
  END r0_rd_out[378]
  PIN r0_rd_out[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 748.945 1511.860 749.015 1512.000 ;
    END
  END r0_rd_out[379]
  PIN r0_rd_out[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 755.025 1511.860 755.095 1512.000 ;
    END
  END r0_rd_out[380]
  PIN r0_rd_out[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 761.105 1511.860 761.175 1512.000 ;
    END
  END r0_rd_out[381]
  PIN r0_rd_out[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 767.185 1511.860 767.255 1512.000 ;
    END
  END r0_rd_out[382]
  PIN r0_rd_out[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 773.265 1511.860 773.335 1512.000 ;
    END
  END r0_rd_out[383]
  PIN r0_rd_out[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 779.345 1511.860 779.415 1512.000 ;
    END
  END r0_rd_out[384]
  PIN r0_rd_out[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 785.425 1511.860 785.495 1512.000 ;
    END
  END r0_rd_out[385]
  PIN r0_rd_out[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 791.505 1511.860 791.575 1512.000 ;
    END
  END r0_rd_out[386]
  PIN r0_rd_out[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 797.585 1511.860 797.655 1512.000 ;
    END
  END r0_rd_out[387]
  PIN r0_rd_out[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 803.665 1511.860 803.735 1512.000 ;
    END
  END r0_rd_out[388]
  PIN r0_rd_out[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 809.745 1511.860 809.815 1512.000 ;
    END
  END r0_rd_out[389]
  PIN r0_rd_out[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 815.825 1511.860 815.895 1512.000 ;
    END
  END r0_rd_out[390]
  PIN r0_rd_out[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 821.905 1511.860 821.975 1512.000 ;
    END
  END r0_rd_out[391]
  PIN r0_rd_out[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 827.985 1511.860 828.055 1512.000 ;
    END
  END r0_rd_out[392]
  PIN r0_rd_out[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 834.065 1511.860 834.135 1512.000 ;
    END
  END r0_rd_out[393]
  PIN r0_rd_out[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 840.145 1511.860 840.215 1512.000 ;
    END
  END r0_rd_out[394]
  PIN r0_rd_out[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 846.225 1511.860 846.295 1512.000 ;
    END
  END r0_rd_out[395]
  PIN r0_rd_out[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 852.305 1511.860 852.375 1512.000 ;
    END
  END r0_rd_out[396]
  PIN r0_rd_out[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 858.385 1511.860 858.455 1512.000 ;
    END
  END r0_rd_out[397]
  PIN r0_rd_out[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 864.465 1511.860 864.535 1512.000 ;
    END
  END r0_rd_out[398]
  PIN r0_rd_out[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 870.545 1511.860 870.615 1512.000 ;
    END
  END r0_rd_out[399]
  PIN r0_rd_out[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 876.625 1511.860 876.695 1512.000 ;
    END
  END r0_rd_out[400]
  PIN r0_rd_out[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 882.705 1511.860 882.775 1512.000 ;
    END
  END r0_rd_out[401]
  PIN r0_rd_out[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 888.785 1511.860 888.855 1512.000 ;
    END
  END r0_rd_out[402]
  PIN r0_rd_out[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 894.865 1511.860 894.935 1512.000 ;
    END
  END r0_rd_out[403]
  PIN r0_rd_out[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 900.945 1511.860 901.015 1512.000 ;
    END
  END r0_rd_out[404]
  PIN r0_rd_out[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 907.025 1511.860 907.095 1512.000 ;
    END
  END r0_rd_out[405]
  PIN r0_rd_out[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 913.105 1511.860 913.175 1512.000 ;
    END
  END r0_rd_out[406]
  PIN r0_rd_out[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 919.185 1511.860 919.255 1512.000 ;
    END
  END r0_rd_out[407]
  PIN r0_rd_out[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 925.265 1511.860 925.335 1512.000 ;
    END
  END r0_rd_out[408]
  PIN r0_rd_out[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 931.345 1511.860 931.415 1512.000 ;
    END
  END r0_rd_out[409]
  PIN r0_rd_out[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 937.425 1511.860 937.495 1512.000 ;
    END
  END r0_rd_out[410]
  PIN r0_rd_out[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 943.505 1511.860 943.575 1512.000 ;
    END
  END r0_rd_out[411]
  PIN r0_rd_out[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 949.585 1511.860 949.655 1512.000 ;
    END
  END r0_rd_out[412]
  PIN r0_rd_out[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 955.665 1511.860 955.735 1512.000 ;
    END
  END r0_rd_out[413]
  PIN r0_rd_out[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 961.745 1511.860 961.815 1512.000 ;
    END
  END r0_rd_out[414]
  PIN r0_rd_out[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 967.825 1511.860 967.895 1512.000 ;
    END
  END r0_rd_out[415]
  PIN r0_rd_out[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 973.905 1511.860 973.975 1512.000 ;
    END
  END r0_rd_out[416]
  PIN r0_rd_out[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 979.985 1511.860 980.055 1512.000 ;
    END
  END r0_rd_out[417]
  PIN r0_rd_out[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 986.065 1511.860 986.135 1512.000 ;
    END
  END r0_rd_out[418]
  PIN r0_rd_out[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 992.145 1511.860 992.215 1512.000 ;
    END
  END r0_rd_out[419]
  PIN r0_rd_out[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 998.225 1511.860 998.295 1512.000 ;
    END
  END r0_rd_out[420]
  PIN r0_rd_out[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1004.305 1511.860 1004.375 1512.000 ;
    END
  END r0_rd_out[421]
  PIN r0_rd_out[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1010.385 1511.860 1010.455 1512.000 ;
    END
  END r0_rd_out[422]
  PIN r0_rd_out[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1016.465 1511.860 1016.535 1512.000 ;
    END
  END r0_rd_out[423]
  PIN r0_rd_out[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1022.545 1511.860 1022.615 1512.000 ;
    END
  END r0_rd_out[424]
  PIN r0_rd_out[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1028.625 1511.860 1028.695 1512.000 ;
    END
  END r0_rd_out[425]
  PIN r0_rd_out[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1034.705 1511.860 1034.775 1512.000 ;
    END
  END r0_rd_out[426]
  PIN r0_rd_out[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1040.785 1511.860 1040.855 1512.000 ;
    END
  END r0_rd_out[427]
  PIN r0_rd_out[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1046.865 1511.860 1046.935 1512.000 ;
    END
  END r0_rd_out[428]
  PIN r0_rd_out[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1052.945 1511.860 1053.015 1512.000 ;
    END
  END r0_rd_out[429]
  PIN r0_rd_out[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1059.025 1511.860 1059.095 1512.000 ;
    END
  END r0_rd_out[430]
  PIN r0_rd_out[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1065.105 1511.860 1065.175 1512.000 ;
    END
  END r0_rd_out[431]
  PIN r0_rd_out[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1071.185 1511.860 1071.255 1512.000 ;
    END
  END r0_rd_out[432]
  PIN r0_rd_out[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1077.265 1511.860 1077.335 1512.000 ;
    END
  END r0_rd_out[433]
  PIN r0_rd_out[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1083.345 1511.860 1083.415 1512.000 ;
    END
  END r0_rd_out[434]
  PIN r0_rd_out[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1089.425 1511.860 1089.495 1512.000 ;
    END
  END r0_rd_out[435]
  PIN r0_rd_out[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1095.505 1511.860 1095.575 1512.000 ;
    END
  END r0_rd_out[436]
  PIN r0_rd_out[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1101.585 1511.860 1101.655 1512.000 ;
    END
  END r0_rd_out[437]
  PIN r0_rd_out[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1107.665 1511.860 1107.735 1512.000 ;
    END
  END r0_rd_out[438]
  PIN r0_rd_out[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1113.745 1511.860 1113.815 1512.000 ;
    END
  END r0_rd_out[439]
  PIN r0_rd_out[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1119.825 1511.860 1119.895 1512.000 ;
    END
  END r0_rd_out[440]
  PIN r0_rd_out[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1125.905 1511.860 1125.975 1512.000 ;
    END
  END r0_rd_out[441]
  PIN r0_rd_out[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1131.985 1511.860 1132.055 1512.000 ;
    END
  END r0_rd_out[442]
  PIN r0_rd_out[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1138.065 1511.860 1138.135 1512.000 ;
    END
  END r0_rd_out[443]
  PIN r0_rd_out[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1144.145 1511.860 1144.215 1512.000 ;
    END
  END r0_rd_out[444]
  PIN r0_rd_out[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1150.225 1511.860 1150.295 1512.000 ;
    END
  END r0_rd_out[445]
  PIN r0_rd_out[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1156.305 1511.860 1156.375 1512.000 ;
    END
  END r0_rd_out[446]
  PIN r0_rd_out[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1162.385 1511.860 1162.455 1512.000 ;
    END
  END r0_rd_out[447]
  PIN r0_rd_out[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1168.465 1511.860 1168.535 1512.000 ;
    END
  END r0_rd_out[448]
  PIN r0_rd_out[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1174.545 1511.860 1174.615 1512.000 ;
    END
  END r0_rd_out[449]
  PIN r0_rd_out[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1180.625 1511.860 1180.695 1512.000 ;
    END
  END r0_rd_out[450]
  PIN r0_rd_out[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1186.705 1511.860 1186.775 1512.000 ;
    END
  END r0_rd_out[451]
  PIN r0_rd_out[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1192.785 1511.860 1192.855 1512.000 ;
    END
  END r0_rd_out[452]
  PIN r0_rd_out[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1198.865 1511.860 1198.935 1512.000 ;
    END
  END r0_rd_out[453]
  PIN r0_rd_out[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1204.945 1511.860 1205.015 1512.000 ;
    END
  END r0_rd_out[454]
  PIN r0_rd_out[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1211.025 1511.860 1211.095 1512.000 ;
    END
  END r0_rd_out[455]
  PIN r0_rd_out[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1217.105 1511.860 1217.175 1512.000 ;
    END
  END r0_rd_out[456]
  PIN r0_rd_out[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1223.185 1511.860 1223.255 1512.000 ;
    END
  END r0_rd_out[457]
  PIN r0_rd_out[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1229.265 1511.860 1229.335 1512.000 ;
    END
  END r0_rd_out[458]
  PIN r0_rd_out[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1235.345 1511.860 1235.415 1512.000 ;
    END
  END r0_rd_out[459]
  PIN r0_rd_out[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1241.425 1511.860 1241.495 1512.000 ;
    END
  END r0_rd_out[460]
  PIN r0_rd_out[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1247.505 1511.860 1247.575 1512.000 ;
    END
  END r0_rd_out[461]
  PIN r0_rd_out[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1253.585 1511.860 1253.655 1512.000 ;
    END
  END r0_rd_out[462]
  PIN r0_rd_out[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1259.665 1511.860 1259.735 1512.000 ;
    END
  END r0_rd_out[463]
  PIN r0_rd_out[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1265.745 1511.860 1265.815 1512.000 ;
    END
  END r0_rd_out[464]
  PIN r0_rd_out[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1271.825 1511.860 1271.895 1512.000 ;
    END
  END r0_rd_out[465]
  PIN r0_rd_out[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1277.905 1511.860 1277.975 1512.000 ;
    END
  END r0_rd_out[466]
  PIN r0_rd_out[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1283.985 1511.860 1284.055 1512.000 ;
    END
  END r0_rd_out[467]
  PIN r0_rd_out[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1290.065 1511.860 1290.135 1512.000 ;
    END
  END r0_rd_out[468]
  PIN r0_rd_out[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1296.145 1511.860 1296.215 1512.000 ;
    END
  END r0_rd_out[469]
  PIN r0_rd_out[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1302.225 1511.860 1302.295 1512.000 ;
    END
  END r0_rd_out[470]
  PIN r0_rd_out[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1308.305 1511.860 1308.375 1512.000 ;
    END
  END r0_rd_out[471]
  PIN r0_rd_out[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1314.385 1511.860 1314.455 1512.000 ;
    END
  END r0_rd_out[472]
  PIN r0_rd_out[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1320.465 1511.860 1320.535 1512.000 ;
    END
  END r0_rd_out[473]
  PIN r0_rd_out[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1326.545 1511.860 1326.615 1512.000 ;
    END
  END r0_rd_out[474]
  PIN r0_rd_out[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1332.625 1511.860 1332.695 1512.000 ;
    END
  END r0_rd_out[475]
  PIN r0_rd_out[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1338.705 1511.860 1338.775 1512.000 ;
    END
  END r0_rd_out[476]
  PIN r0_rd_out[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1344.785 1511.860 1344.855 1512.000 ;
    END
  END r0_rd_out[477]
  PIN r0_rd_out[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1350.865 1511.860 1350.935 1512.000 ;
    END
  END r0_rd_out[478]
  PIN r0_rd_out[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1356.945 1511.860 1357.015 1512.000 ;
    END
  END r0_rd_out[479]
  PIN r0_rd_out[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1363.025 1511.860 1363.095 1512.000 ;
    END
  END r0_rd_out[480]
  PIN r0_rd_out[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1369.105 1511.860 1369.175 1512.000 ;
    END
  END r0_rd_out[481]
  PIN r0_rd_out[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1375.185 1511.860 1375.255 1512.000 ;
    END
  END r0_rd_out[482]
  PIN r0_rd_out[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1381.265 1511.860 1381.335 1512.000 ;
    END
  END r0_rd_out[483]
  PIN r0_rd_out[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1387.345 1511.860 1387.415 1512.000 ;
    END
  END r0_rd_out[484]
  PIN r0_rd_out[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1393.425 1511.860 1393.495 1512.000 ;
    END
  END r0_rd_out[485]
  PIN r0_rd_out[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1399.505 1511.860 1399.575 1512.000 ;
    END
  END r0_rd_out[486]
  PIN r0_rd_out[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1405.585 1511.860 1405.655 1512.000 ;
    END
  END r0_rd_out[487]
  PIN r0_rd_out[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1411.665 1511.860 1411.735 1512.000 ;
    END
  END r0_rd_out[488]
  PIN r0_rd_out[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1417.745 1511.860 1417.815 1512.000 ;
    END
  END r0_rd_out[489]
  PIN r0_rd_out[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1423.825 1511.860 1423.895 1512.000 ;
    END
  END r0_rd_out[490]
  PIN r0_rd_out[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1429.905 1511.860 1429.975 1512.000 ;
    END
  END r0_rd_out[491]
  PIN r0_rd_out[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1435.985 1511.860 1436.055 1512.000 ;
    END
  END r0_rd_out[492]
  PIN r0_rd_out[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1442.065 1511.860 1442.135 1512.000 ;
    END
  END r0_rd_out[493]
  PIN r0_rd_out[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1448.145 1511.860 1448.215 1512.000 ;
    END
  END r0_rd_out[494]
  PIN r0_rd_out[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1454.225 1511.860 1454.295 1512.000 ;
    END
  END r0_rd_out[495]
  PIN r0_rd_out[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1460.305 1511.860 1460.375 1512.000 ;
    END
  END r0_rd_out[496]
  PIN r0_rd_out[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1466.385 1511.860 1466.455 1512.000 ;
    END
  END r0_rd_out[497]
  PIN r0_rd_out[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1472.465 1511.860 1472.535 1512.000 ;
    END
  END r0_rd_out[498]
  PIN r0_rd_out[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1478.545 1511.860 1478.615 1512.000 ;
    END
  END r0_rd_out[499]
  PIN r0_rd_out[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1484.625 1511.860 1484.695 1512.000 ;
    END
  END r0_rd_out[500]
  PIN r0_rd_out[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1490.705 1511.860 1490.775 1512.000 ;
    END
  END r0_rd_out[501]
  PIN r0_rd_out[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1496.785 1511.860 1496.855 1512.000 ;
    END
  END r0_rd_out[502]
  PIN r0_rd_out[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1502.865 1511.860 1502.935 1512.000 ;
    END
  END r0_rd_out[503]
  PIN r0_rd_out[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1508.945 1511.860 1509.015 1512.000 ;
    END
  END r0_rd_out[504]
  PIN r0_rd_out[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1515.025 1511.860 1515.095 1512.000 ;
    END
  END r0_rd_out[505]
  PIN r0_rd_out[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1521.105 1511.860 1521.175 1512.000 ;
    END
  END r0_rd_out[506]
  PIN r0_rd_out[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1527.185 1511.860 1527.255 1512.000 ;
    END
  END r0_rd_out[507]
  PIN r0_rd_out[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1533.265 1511.860 1533.335 1512.000 ;
    END
  END r0_rd_out[508]
  PIN r0_rd_out[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1539.345 1511.860 1539.415 1512.000 ;
    END
  END r0_rd_out[509]
  PIN r0_rd_out[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1545.425 1511.860 1545.495 1512.000 ;
    END
  END r0_rd_out[510]
  PIN r0_rd_out[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1551.505 1511.860 1551.575 1512.000 ;
    END
  END r0_rd_out[511]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1380.645 0.140 1380.715 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1391.425 0.140 1391.495 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1402.205 0.140 1402.275 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1412.985 0.140 1413.055 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1423.765 0.140 1423.835 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1434.545 0.140 1434.615 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1380.645 1609.300 1380.715 ;
    END
  END w0_addr_in[6]
  PIN w0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1391.425 1609.300 1391.495 ;
    END
  END w0_addr_in[7]
  PIN w0_addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1402.205 1609.300 1402.275 ;
    END
  END w0_addr_in[8]
  PIN w0_addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1412.985 1609.300 1413.055 ;
    END
  END w0_addr_in[9]
  PIN w0_addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1423.765 1609.300 1423.835 ;
    END
  END w0_addr_in[10]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1445.325 0.140 1445.395 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1456.105 0.140 1456.175 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1466.885 0.140 1466.955 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1477.665 0.140 1477.735 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1488.445 0.140 1488.515 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1499.225 0.140 1499.295 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1434.545 1609.300 1434.615 ;
    END
  END r0_addr_in[6]
  PIN r0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1445.325 1609.300 1445.395 ;
    END
  END r0_addr_in[7]
  PIN r0_addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1456.105 1609.300 1456.175 ;
    END
  END r0_addr_in[8]
  PIN r0_addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1466.885 1609.300 1466.955 ;
    END
  END r0_addr_in[9]
  PIN r0_addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 1609.160 1477.665 1609.300 1477.735 ;
    END
  END r0_addr_in[10]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1557.585 1511.860 1557.655 1512.000 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1563.665 1511.860 1563.735 1512.000 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1569.745 1511.860 1569.815 1512.000 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1575.825 1511.860 1575.895 1512.000 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
      RECT 1581.905 1511.860 1581.975 1512.000 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 0.430 0.700 0.710 1511.300 ;
      RECT 2.670 0.700 2.950 1511.300 ;
      RECT 4.910 0.700 5.190 1511.300 ;
      RECT 7.150 0.700 7.430 1511.300 ;
      RECT 9.390 0.700 9.670 1511.300 ;
      RECT 11.630 0.700 11.910 1511.300 ;
      RECT 13.870 0.700 14.150 1511.300 ;
      RECT 16.110 0.700 16.390 1511.300 ;
      RECT 18.350 0.700 18.630 1511.300 ;
      RECT 20.590 0.700 20.870 1511.300 ;
      RECT 22.830 0.700 23.110 1511.300 ;
      RECT 25.070 0.700 25.350 1511.300 ;
      RECT 27.310 0.700 27.590 1511.300 ;
      RECT 29.550 0.700 29.830 1511.300 ;
      RECT 31.790 0.700 32.070 1511.300 ;
      RECT 34.030 0.700 34.310 1511.300 ;
      RECT 36.270 0.700 36.550 1511.300 ;
      RECT 38.510 0.700 38.790 1511.300 ;
      RECT 40.750 0.700 41.030 1511.300 ;
      RECT 42.990 0.700 43.270 1511.300 ;
      RECT 45.230 0.700 45.510 1511.300 ;
      RECT 47.470 0.700 47.750 1511.300 ;
      RECT 49.710 0.700 49.990 1511.300 ;
      RECT 51.950 0.700 52.230 1511.300 ;
      RECT 54.190 0.700 54.470 1511.300 ;
      RECT 56.430 0.700 56.710 1511.300 ;
      RECT 58.670 0.700 58.950 1511.300 ;
      RECT 60.910 0.700 61.190 1511.300 ;
      RECT 63.150 0.700 63.430 1511.300 ;
      RECT 65.390 0.700 65.670 1511.300 ;
      RECT 67.630 0.700 67.910 1511.300 ;
      RECT 69.870 0.700 70.150 1511.300 ;
      RECT 72.110 0.700 72.390 1511.300 ;
      RECT 74.350 0.700 74.630 1511.300 ;
      RECT 76.590 0.700 76.870 1511.300 ;
      RECT 78.830 0.700 79.110 1511.300 ;
      RECT 81.070 0.700 81.350 1511.300 ;
      RECT 83.310 0.700 83.590 1511.300 ;
      RECT 85.550 0.700 85.830 1511.300 ;
      RECT 87.790 0.700 88.070 1511.300 ;
      RECT 90.030 0.700 90.310 1511.300 ;
      RECT 92.270 0.700 92.550 1511.300 ;
      RECT 94.510 0.700 94.790 1511.300 ;
      RECT 96.750 0.700 97.030 1511.300 ;
      RECT 98.990 0.700 99.270 1511.300 ;
      RECT 101.230 0.700 101.510 1511.300 ;
      RECT 103.470 0.700 103.750 1511.300 ;
      RECT 105.710 0.700 105.990 1511.300 ;
      RECT 107.950 0.700 108.230 1511.300 ;
      RECT 110.190 0.700 110.470 1511.300 ;
      RECT 112.430 0.700 112.710 1511.300 ;
      RECT 114.670 0.700 114.950 1511.300 ;
      RECT 116.910 0.700 117.190 1511.300 ;
      RECT 119.150 0.700 119.430 1511.300 ;
      RECT 121.390 0.700 121.670 1511.300 ;
      RECT 123.630 0.700 123.910 1511.300 ;
      RECT 125.870 0.700 126.150 1511.300 ;
      RECT 128.110 0.700 128.390 1511.300 ;
      RECT 130.350 0.700 130.630 1511.300 ;
      RECT 132.590 0.700 132.870 1511.300 ;
      RECT 134.830 0.700 135.110 1511.300 ;
      RECT 137.070 0.700 137.350 1511.300 ;
      RECT 139.310 0.700 139.590 1511.300 ;
      RECT 141.550 0.700 141.830 1511.300 ;
      RECT 143.790 0.700 144.070 1511.300 ;
      RECT 146.030 0.700 146.310 1511.300 ;
      RECT 148.270 0.700 148.550 1511.300 ;
      RECT 150.510 0.700 150.790 1511.300 ;
      RECT 152.750 0.700 153.030 1511.300 ;
      RECT 154.990 0.700 155.270 1511.300 ;
      RECT 157.230 0.700 157.510 1511.300 ;
      RECT 159.470 0.700 159.750 1511.300 ;
      RECT 161.710 0.700 161.990 1511.300 ;
      RECT 163.950 0.700 164.230 1511.300 ;
      RECT 166.190 0.700 166.470 1511.300 ;
      RECT 168.430 0.700 168.710 1511.300 ;
      RECT 170.670 0.700 170.950 1511.300 ;
      RECT 172.910 0.700 173.190 1511.300 ;
      RECT 175.150 0.700 175.430 1511.300 ;
      RECT 177.390 0.700 177.670 1511.300 ;
      RECT 179.630 0.700 179.910 1511.300 ;
      RECT 181.870 0.700 182.150 1511.300 ;
      RECT 184.110 0.700 184.390 1511.300 ;
      RECT 186.350 0.700 186.630 1511.300 ;
      RECT 188.590 0.700 188.870 1511.300 ;
      RECT 190.830 0.700 191.110 1511.300 ;
      RECT 193.070 0.700 193.350 1511.300 ;
      RECT 195.310 0.700 195.590 1511.300 ;
      RECT 197.550 0.700 197.830 1511.300 ;
      RECT 199.790 0.700 200.070 1511.300 ;
      RECT 202.030 0.700 202.310 1511.300 ;
      RECT 204.270 0.700 204.550 1511.300 ;
      RECT 206.510 0.700 206.790 1511.300 ;
      RECT 208.750 0.700 209.030 1511.300 ;
      RECT 210.990 0.700 211.270 1511.300 ;
      RECT 213.230 0.700 213.510 1511.300 ;
      RECT 215.470 0.700 215.750 1511.300 ;
      RECT 217.710 0.700 217.990 1511.300 ;
      RECT 219.950 0.700 220.230 1511.300 ;
      RECT 222.190 0.700 222.470 1511.300 ;
      RECT 224.430 0.700 224.710 1511.300 ;
      RECT 226.670 0.700 226.950 1511.300 ;
      RECT 228.910 0.700 229.190 1511.300 ;
      RECT 231.150 0.700 231.430 1511.300 ;
      RECT 233.390 0.700 233.670 1511.300 ;
      RECT 235.630 0.700 235.910 1511.300 ;
      RECT 237.870 0.700 238.150 1511.300 ;
      RECT 240.110 0.700 240.390 1511.300 ;
      RECT 242.350 0.700 242.630 1511.300 ;
      RECT 244.590 0.700 244.870 1511.300 ;
      RECT 246.830 0.700 247.110 1511.300 ;
      RECT 249.070 0.700 249.350 1511.300 ;
      RECT 251.310 0.700 251.590 1511.300 ;
      RECT 253.550 0.700 253.830 1511.300 ;
      RECT 255.790 0.700 256.070 1511.300 ;
      RECT 258.030 0.700 258.310 1511.300 ;
      RECT 260.270 0.700 260.550 1511.300 ;
      RECT 262.510 0.700 262.790 1511.300 ;
      RECT 264.750 0.700 265.030 1511.300 ;
      RECT 266.990 0.700 267.270 1511.300 ;
      RECT 269.230 0.700 269.510 1511.300 ;
      RECT 271.470 0.700 271.750 1511.300 ;
      RECT 273.710 0.700 273.990 1511.300 ;
      RECT 275.950 0.700 276.230 1511.300 ;
      RECT 278.190 0.700 278.470 1511.300 ;
      RECT 280.430 0.700 280.710 1511.300 ;
      RECT 282.670 0.700 282.950 1511.300 ;
      RECT 284.910 0.700 285.190 1511.300 ;
      RECT 287.150 0.700 287.430 1511.300 ;
      RECT 289.390 0.700 289.670 1511.300 ;
      RECT 291.630 0.700 291.910 1511.300 ;
      RECT 293.870 0.700 294.150 1511.300 ;
      RECT 296.110 0.700 296.390 1511.300 ;
      RECT 298.350 0.700 298.630 1511.300 ;
      RECT 300.590 0.700 300.870 1511.300 ;
      RECT 302.830 0.700 303.110 1511.300 ;
      RECT 305.070 0.700 305.350 1511.300 ;
      RECT 307.310 0.700 307.590 1511.300 ;
      RECT 309.550 0.700 309.830 1511.300 ;
      RECT 311.790 0.700 312.070 1511.300 ;
      RECT 314.030 0.700 314.310 1511.300 ;
      RECT 316.270 0.700 316.550 1511.300 ;
      RECT 318.510 0.700 318.790 1511.300 ;
      RECT 320.750 0.700 321.030 1511.300 ;
      RECT 322.990 0.700 323.270 1511.300 ;
      RECT 325.230 0.700 325.510 1511.300 ;
      RECT 327.470 0.700 327.750 1511.300 ;
      RECT 329.710 0.700 329.990 1511.300 ;
      RECT 331.950 0.700 332.230 1511.300 ;
      RECT 334.190 0.700 334.470 1511.300 ;
      RECT 336.430 0.700 336.710 1511.300 ;
      RECT 338.670 0.700 338.950 1511.300 ;
      RECT 340.910 0.700 341.190 1511.300 ;
      RECT 343.150 0.700 343.430 1511.300 ;
      RECT 345.390 0.700 345.670 1511.300 ;
      RECT 347.630 0.700 347.910 1511.300 ;
      RECT 349.870 0.700 350.150 1511.300 ;
      RECT 352.110 0.700 352.390 1511.300 ;
      RECT 354.350 0.700 354.630 1511.300 ;
      RECT 356.590 0.700 356.870 1511.300 ;
      RECT 358.830 0.700 359.110 1511.300 ;
      RECT 361.070 0.700 361.350 1511.300 ;
      RECT 363.310 0.700 363.590 1511.300 ;
      RECT 365.550 0.700 365.830 1511.300 ;
      RECT 367.790 0.700 368.070 1511.300 ;
      RECT 370.030 0.700 370.310 1511.300 ;
      RECT 372.270 0.700 372.550 1511.300 ;
      RECT 374.510 0.700 374.790 1511.300 ;
      RECT 376.750 0.700 377.030 1511.300 ;
      RECT 378.990 0.700 379.270 1511.300 ;
      RECT 381.230 0.700 381.510 1511.300 ;
      RECT 383.470 0.700 383.750 1511.300 ;
      RECT 385.710 0.700 385.990 1511.300 ;
      RECT 387.950 0.700 388.230 1511.300 ;
      RECT 390.190 0.700 390.470 1511.300 ;
      RECT 392.430 0.700 392.710 1511.300 ;
      RECT 394.670 0.700 394.950 1511.300 ;
      RECT 396.910 0.700 397.190 1511.300 ;
      RECT 399.150 0.700 399.430 1511.300 ;
      RECT 401.390 0.700 401.670 1511.300 ;
      RECT 403.630 0.700 403.910 1511.300 ;
      RECT 405.870 0.700 406.150 1511.300 ;
      RECT 408.110 0.700 408.390 1511.300 ;
      RECT 410.350 0.700 410.630 1511.300 ;
      RECT 412.590 0.700 412.870 1511.300 ;
      RECT 414.830 0.700 415.110 1511.300 ;
      RECT 417.070 0.700 417.350 1511.300 ;
      RECT 419.310 0.700 419.590 1511.300 ;
      RECT 421.550 0.700 421.830 1511.300 ;
      RECT 423.790 0.700 424.070 1511.300 ;
      RECT 426.030 0.700 426.310 1511.300 ;
      RECT 428.270 0.700 428.550 1511.300 ;
      RECT 430.510 0.700 430.790 1511.300 ;
      RECT 432.750 0.700 433.030 1511.300 ;
      RECT 434.990 0.700 435.270 1511.300 ;
      RECT 437.230 0.700 437.510 1511.300 ;
      RECT 439.470 0.700 439.750 1511.300 ;
      RECT 441.710 0.700 441.990 1511.300 ;
      RECT 443.950 0.700 444.230 1511.300 ;
      RECT 446.190 0.700 446.470 1511.300 ;
      RECT 448.430 0.700 448.710 1511.300 ;
      RECT 450.670 0.700 450.950 1511.300 ;
      RECT 452.910 0.700 453.190 1511.300 ;
      RECT 455.150 0.700 455.430 1511.300 ;
      RECT 457.390 0.700 457.670 1511.300 ;
      RECT 459.630 0.700 459.910 1511.300 ;
      RECT 461.870 0.700 462.150 1511.300 ;
      RECT 464.110 0.700 464.390 1511.300 ;
      RECT 466.350 0.700 466.630 1511.300 ;
      RECT 468.590 0.700 468.870 1511.300 ;
      RECT 470.830 0.700 471.110 1511.300 ;
      RECT 473.070 0.700 473.350 1511.300 ;
      RECT 475.310 0.700 475.590 1511.300 ;
      RECT 477.550 0.700 477.830 1511.300 ;
      RECT 479.790 0.700 480.070 1511.300 ;
      RECT 482.030 0.700 482.310 1511.300 ;
      RECT 484.270 0.700 484.550 1511.300 ;
      RECT 486.510 0.700 486.790 1511.300 ;
      RECT 488.750 0.700 489.030 1511.300 ;
      RECT 490.990 0.700 491.270 1511.300 ;
      RECT 493.230 0.700 493.510 1511.300 ;
      RECT 495.470 0.700 495.750 1511.300 ;
      RECT 497.710 0.700 497.990 1511.300 ;
      RECT 499.950 0.700 500.230 1511.300 ;
      RECT 502.190 0.700 502.470 1511.300 ;
      RECT 504.430 0.700 504.710 1511.300 ;
      RECT 506.670 0.700 506.950 1511.300 ;
      RECT 508.910 0.700 509.190 1511.300 ;
      RECT 511.150 0.700 511.430 1511.300 ;
      RECT 513.390 0.700 513.670 1511.300 ;
      RECT 515.630 0.700 515.910 1511.300 ;
      RECT 517.870 0.700 518.150 1511.300 ;
      RECT 520.110 0.700 520.390 1511.300 ;
      RECT 522.350 0.700 522.630 1511.300 ;
      RECT 524.590 0.700 524.870 1511.300 ;
      RECT 526.830 0.700 527.110 1511.300 ;
      RECT 529.070 0.700 529.350 1511.300 ;
      RECT 531.310 0.700 531.590 1511.300 ;
      RECT 533.550 0.700 533.830 1511.300 ;
      RECT 535.790 0.700 536.070 1511.300 ;
      RECT 538.030 0.700 538.310 1511.300 ;
      RECT 540.270 0.700 540.550 1511.300 ;
      RECT 542.510 0.700 542.790 1511.300 ;
      RECT 544.750 0.700 545.030 1511.300 ;
      RECT 546.990 0.700 547.270 1511.300 ;
      RECT 549.230 0.700 549.510 1511.300 ;
      RECT 551.470 0.700 551.750 1511.300 ;
      RECT 553.710 0.700 553.990 1511.300 ;
      RECT 555.950 0.700 556.230 1511.300 ;
      RECT 558.190 0.700 558.470 1511.300 ;
      RECT 560.430 0.700 560.710 1511.300 ;
      RECT 562.670 0.700 562.950 1511.300 ;
      RECT 564.910 0.700 565.190 1511.300 ;
      RECT 567.150 0.700 567.430 1511.300 ;
      RECT 569.390 0.700 569.670 1511.300 ;
      RECT 571.630 0.700 571.910 1511.300 ;
      RECT 573.870 0.700 574.150 1511.300 ;
      RECT 576.110 0.700 576.390 1511.300 ;
      RECT 578.350 0.700 578.630 1511.300 ;
      RECT 580.590 0.700 580.870 1511.300 ;
      RECT 582.830 0.700 583.110 1511.300 ;
      RECT 585.070 0.700 585.350 1511.300 ;
      RECT 587.310 0.700 587.590 1511.300 ;
      RECT 589.550 0.700 589.830 1511.300 ;
      RECT 591.790 0.700 592.070 1511.300 ;
      RECT 594.030 0.700 594.310 1511.300 ;
      RECT 596.270 0.700 596.550 1511.300 ;
      RECT 598.510 0.700 598.790 1511.300 ;
      RECT 600.750 0.700 601.030 1511.300 ;
      RECT 602.990 0.700 603.270 1511.300 ;
      RECT 605.230 0.700 605.510 1511.300 ;
      RECT 607.470 0.700 607.750 1511.300 ;
      RECT 609.710 0.700 609.990 1511.300 ;
      RECT 611.950 0.700 612.230 1511.300 ;
      RECT 614.190 0.700 614.470 1511.300 ;
      RECT 616.430 0.700 616.710 1511.300 ;
      RECT 618.670 0.700 618.950 1511.300 ;
      RECT 620.910 0.700 621.190 1511.300 ;
      RECT 623.150 0.700 623.430 1511.300 ;
      RECT 625.390 0.700 625.670 1511.300 ;
      RECT 627.630 0.700 627.910 1511.300 ;
      RECT 629.870 0.700 630.150 1511.300 ;
      RECT 632.110 0.700 632.390 1511.300 ;
      RECT 634.350 0.700 634.630 1511.300 ;
      RECT 636.590 0.700 636.870 1511.300 ;
      RECT 638.830 0.700 639.110 1511.300 ;
      RECT 641.070 0.700 641.350 1511.300 ;
      RECT 643.310 0.700 643.590 1511.300 ;
      RECT 645.550 0.700 645.830 1511.300 ;
      RECT 647.790 0.700 648.070 1511.300 ;
      RECT 650.030 0.700 650.310 1511.300 ;
      RECT 652.270 0.700 652.550 1511.300 ;
      RECT 654.510 0.700 654.790 1511.300 ;
      RECT 656.750 0.700 657.030 1511.300 ;
      RECT 658.990 0.700 659.270 1511.300 ;
      RECT 661.230 0.700 661.510 1511.300 ;
      RECT 663.470 0.700 663.750 1511.300 ;
      RECT 665.710 0.700 665.990 1511.300 ;
      RECT 667.950 0.700 668.230 1511.300 ;
      RECT 670.190 0.700 670.470 1511.300 ;
      RECT 672.430 0.700 672.710 1511.300 ;
      RECT 674.670 0.700 674.950 1511.300 ;
      RECT 676.910 0.700 677.190 1511.300 ;
      RECT 679.150 0.700 679.430 1511.300 ;
      RECT 681.390 0.700 681.670 1511.300 ;
      RECT 683.630 0.700 683.910 1511.300 ;
      RECT 685.870 0.700 686.150 1511.300 ;
      RECT 688.110 0.700 688.390 1511.300 ;
      RECT 690.350 0.700 690.630 1511.300 ;
      RECT 692.590 0.700 692.870 1511.300 ;
      RECT 694.830 0.700 695.110 1511.300 ;
      RECT 697.070 0.700 697.350 1511.300 ;
      RECT 699.310 0.700 699.590 1511.300 ;
      RECT 701.550 0.700 701.830 1511.300 ;
      RECT 703.790 0.700 704.070 1511.300 ;
      RECT 706.030 0.700 706.310 1511.300 ;
      RECT 708.270 0.700 708.550 1511.300 ;
      RECT 710.510 0.700 710.790 1511.300 ;
      RECT 712.750 0.700 713.030 1511.300 ;
      RECT 714.990 0.700 715.270 1511.300 ;
      RECT 717.230 0.700 717.510 1511.300 ;
      RECT 719.470 0.700 719.750 1511.300 ;
      RECT 721.710 0.700 721.990 1511.300 ;
      RECT 723.950 0.700 724.230 1511.300 ;
      RECT 726.190 0.700 726.470 1511.300 ;
      RECT 728.430 0.700 728.710 1511.300 ;
      RECT 730.670 0.700 730.950 1511.300 ;
      RECT 732.910 0.700 733.190 1511.300 ;
      RECT 735.150 0.700 735.430 1511.300 ;
      RECT 737.390 0.700 737.670 1511.300 ;
      RECT 739.630 0.700 739.910 1511.300 ;
      RECT 741.870 0.700 742.150 1511.300 ;
      RECT 744.110 0.700 744.390 1511.300 ;
      RECT 746.350 0.700 746.630 1511.300 ;
      RECT 748.590 0.700 748.870 1511.300 ;
      RECT 750.830 0.700 751.110 1511.300 ;
      RECT 753.070 0.700 753.350 1511.300 ;
      RECT 755.310 0.700 755.590 1511.300 ;
      RECT 757.550 0.700 757.830 1511.300 ;
      RECT 759.790 0.700 760.070 1511.300 ;
      RECT 762.030 0.700 762.310 1511.300 ;
      RECT 764.270 0.700 764.550 1511.300 ;
      RECT 766.510 0.700 766.790 1511.300 ;
      RECT 768.750 0.700 769.030 1511.300 ;
      RECT 770.990 0.700 771.270 1511.300 ;
      RECT 773.230 0.700 773.510 1511.300 ;
      RECT 775.470 0.700 775.750 1511.300 ;
      RECT 777.710 0.700 777.990 1511.300 ;
      RECT 779.950 0.700 780.230 1511.300 ;
      RECT 782.190 0.700 782.470 1511.300 ;
      RECT 784.430 0.700 784.710 1511.300 ;
      RECT 786.670 0.700 786.950 1511.300 ;
      RECT 788.910 0.700 789.190 1511.300 ;
      RECT 791.150 0.700 791.430 1511.300 ;
      RECT 793.390 0.700 793.670 1511.300 ;
      RECT 795.630 0.700 795.910 1511.300 ;
      RECT 797.870 0.700 798.150 1511.300 ;
      RECT 800.110 0.700 800.390 1511.300 ;
      RECT 802.350 0.700 802.630 1511.300 ;
      RECT 804.590 0.700 804.870 1511.300 ;
      RECT 806.830 0.700 807.110 1511.300 ;
      RECT 809.070 0.700 809.350 1511.300 ;
      RECT 811.310 0.700 811.590 1511.300 ;
      RECT 813.550 0.700 813.830 1511.300 ;
      RECT 815.790 0.700 816.070 1511.300 ;
      RECT 818.030 0.700 818.310 1511.300 ;
      RECT 820.270 0.700 820.550 1511.300 ;
      RECT 822.510 0.700 822.790 1511.300 ;
      RECT 824.750 0.700 825.030 1511.300 ;
      RECT 826.990 0.700 827.270 1511.300 ;
      RECT 829.230 0.700 829.510 1511.300 ;
      RECT 831.470 0.700 831.750 1511.300 ;
      RECT 833.710 0.700 833.990 1511.300 ;
      RECT 835.950 0.700 836.230 1511.300 ;
      RECT 838.190 0.700 838.470 1511.300 ;
      RECT 840.430 0.700 840.710 1511.300 ;
      RECT 842.670 0.700 842.950 1511.300 ;
      RECT 844.910 0.700 845.190 1511.300 ;
      RECT 847.150 0.700 847.430 1511.300 ;
      RECT 849.390 0.700 849.670 1511.300 ;
      RECT 851.630 0.700 851.910 1511.300 ;
      RECT 853.870 0.700 854.150 1511.300 ;
      RECT 856.110 0.700 856.390 1511.300 ;
      RECT 858.350 0.700 858.630 1511.300 ;
      RECT 860.590 0.700 860.870 1511.300 ;
      RECT 862.830 0.700 863.110 1511.300 ;
      RECT 865.070 0.700 865.350 1511.300 ;
      RECT 867.310 0.700 867.590 1511.300 ;
      RECT 869.550 0.700 869.830 1511.300 ;
      RECT 871.790 0.700 872.070 1511.300 ;
      RECT 874.030 0.700 874.310 1511.300 ;
      RECT 876.270 0.700 876.550 1511.300 ;
      RECT 878.510 0.700 878.790 1511.300 ;
      RECT 880.750 0.700 881.030 1511.300 ;
      RECT 882.990 0.700 883.270 1511.300 ;
      RECT 885.230 0.700 885.510 1511.300 ;
      RECT 887.470 0.700 887.750 1511.300 ;
      RECT 889.710 0.700 889.990 1511.300 ;
      RECT 891.950 0.700 892.230 1511.300 ;
      RECT 894.190 0.700 894.470 1511.300 ;
      RECT 896.430 0.700 896.710 1511.300 ;
      RECT 898.670 0.700 898.950 1511.300 ;
      RECT 900.910 0.700 901.190 1511.300 ;
      RECT 903.150 0.700 903.430 1511.300 ;
      RECT 905.390 0.700 905.670 1511.300 ;
      RECT 907.630 0.700 907.910 1511.300 ;
      RECT 909.870 0.700 910.150 1511.300 ;
      RECT 912.110 0.700 912.390 1511.300 ;
      RECT 914.350 0.700 914.630 1511.300 ;
      RECT 916.590 0.700 916.870 1511.300 ;
      RECT 918.830 0.700 919.110 1511.300 ;
      RECT 921.070 0.700 921.350 1511.300 ;
      RECT 923.310 0.700 923.590 1511.300 ;
      RECT 925.550 0.700 925.830 1511.300 ;
      RECT 927.790 0.700 928.070 1511.300 ;
      RECT 930.030 0.700 930.310 1511.300 ;
      RECT 932.270 0.700 932.550 1511.300 ;
      RECT 934.510 0.700 934.790 1511.300 ;
      RECT 936.750 0.700 937.030 1511.300 ;
      RECT 938.990 0.700 939.270 1511.300 ;
      RECT 941.230 0.700 941.510 1511.300 ;
      RECT 943.470 0.700 943.750 1511.300 ;
      RECT 945.710 0.700 945.990 1511.300 ;
      RECT 947.950 0.700 948.230 1511.300 ;
      RECT 950.190 0.700 950.470 1511.300 ;
      RECT 952.430 0.700 952.710 1511.300 ;
      RECT 954.670 0.700 954.950 1511.300 ;
      RECT 956.910 0.700 957.190 1511.300 ;
      RECT 959.150 0.700 959.430 1511.300 ;
      RECT 961.390 0.700 961.670 1511.300 ;
      RECT 963.630 0.700 963.910 1511.300 ;
      RECT 965.870 0.700 966.150 1511.300 ;
      RECT 968.110 0.700 968.390 1511.300 ;
      RECT 970.350 0.700 970.630 1511.300 ;
      RECT 972.590 0.700 972.870 1511.300 ;
      RECT 974.830 0.700 975.110 1511.300 ;
      RECT 977.070 0.700 977.350 1511.300 ;
      RECT 979.310 0.700 979.590 1511.300 ;
      RECT 981.550 0.700 981.830 1511.300 ;
      RECT 983.790 0.700 984.070 1511.300 ;
      RECT 986.030 0.700 986.310 1511.300 ;
      RECT 988.270 0.700 988.550 1511.300 ;
      RECT 990.510 0.700 990.790 1511.300 ;
      RECT 992.750 0.700 993.030 1511.300 ;
      RECT 994.990 0.700 995.270 1511.300 ;
      RECT 997.230 0.700 997.510 1511.300 ;
      RECT 999.470 0.700 999.750 1511.300 ;
      RECT 1001.710 0.700 1001.990 1511.300 ;
      RECT 1003.950 0.700 1004.230 1511.300 ;
      RECT 1006.190 0.700 1006.470 1511.300 ;
      RECT 1008.430 0.700 1008.710 1511.300 ;
      RECT 1010.670 0.700 1010.950 1511.300 ;
      RECT 1012.910 0.700 1013.190 1511.300 ;
      RECT 1015.150 0.700 1015.430 1511.300 ;
      RECT 1017.390 0.700 1017.670 1511.300 ;
      RECT 1019.630 0.700 1019.910 1511.300 ;
      RECT 1021.870 0.700 1022.150 1511.300 ;
      RECT 1024.110 0.700 1024.390 1511.300 ;
      RECT 1026.350 0.700 1026.630 1511.300 ;
      RECT 1028.590 0.700 1028.870 1511.300 ;
      RECT 1030.830 0.700 1031.110 1511.300 ;
      RECT 1033.070 0.700 1033.350 1511.300 ;
      RECT 1035.310 0.700 1035.590 1511.300 ;
      RECT 1037.550 0.700 1037.830 1511.300 ;
      RECT 1039.790 0.700 1040.070 1511.300 ;
      RECT 1042.030 0.700 1042.310 1511.300 ;
      RECT 1044.270 0.700 1044.550 1511.300 ;
      RECT 1046.510 0.700 1046.790 1511.300 ;
      RECT 1048.750 0.700 1049.030 1511.300 ;
      RECT 1050.990 0.700 1051.270 1511.300 ;
      RECT 1053.230 0.700 1053.510 1511.300 ;
      RECT 1055.470 0.700 1055.750 1511.300 ;
      RECT 1057.710 0.700 1057.990 1511.300 ;
      RECT 1059.950 0.700 1060.230 1511.300 ;
      RECT 1062.190 0.700 1062.470 1511.300 ;
      RECT 1064.430 0.700 1064.710 1511.300 ;
      RECT 1066.670 0.700 1066.950 1511.300 ;
      RECT 1068.910 0.700 1069.190 1511.300 ;
      RECT 1071.150 0.700 1071.430 1511.300 ;
      RECT 1073.390 0.700 1073.670 1511.300 ;
      RECT 1075.630 0.700 1075.910 1511.300 ;
      RECT 1077.870 0.700 1078.150 1511.300 ;
      RECT 1080.110 0.700 1080.390 1511.300 ;
      RECT 1082.350 0.700 1082.630 1511.300 ;
      RECT 1084.590 0.700 1084.870 1511.300 ;
      RECT 1086.830 0.700 1087.110 1511.300 ;
      RECT 1089.070 0.700 1089.350 1511.300 ;
      RECT 1091.310 0.700 1091.590 1511.300 ;
      RECT 1093.550 0.700 1093.830 1511.300 ;
      RECT 1095.790 0.700 1096.070 1511.300 ;
      RECT 1098.030 0.700 1098.310 1511.300 ;
      RECT 1100.270 0.700 1100.550 1511.300 ;
      RECT 1102.510 0.700 1102.790 1511.300 ;
      RECT 1104.750 0.700 1105.030 1511.300 ;
      RECT 1106.990 0.700 1107.270 1511.300 ;
      RECT 1109.230 0.700 1109.510 1511.300 ;
      RECT 1111.470 0.700 1111.750 1511.300 ;
      RECT 1113.710 0.700 1113.990 1511.300 ;
      RECT 1115.950 0.700 1116.230 1511.300 ;
      RECT 1118.190 0.700 1118.470 1511.300 ;
      RECT 1120.430 0.700 1120.710 1511.300 ;
      RECT 1122.670 0.700 1122.950 1511.300 ;
      RECT 1124.910 0.700 1125.190 1511.300 ;
      RECT 1127.150 0.700 1127.430 1511.300 ;
      RECT 1129.390 0.700 1129.670 1511.300 ;
      RECT 1131.630 0.700 1131.910 1511.300 ;
      RECT 1133.870 0.700 1134.150 1511.300 ;
      RECT 1136.110 0.700 1136.390 1511.300 ;
      RECT 1138.350 0.700 1138.630 1511.300 ;
      RECT 1140.590 0.700 1140.870 1511.300 ;
      RECT 1142.830 0.700 1143.110 1511.300 ;
      RECT 1145.070 0.700 1145.350 1511.300 ;
      RECT 1147.310 0.700 1147.590 1511.300 ;
      RECT 1149.550 0.700 1149.830 1511.300 ;
      RECT 1151.790 0.700 1152.070 1511.300 ;
      RECT 1154.030 0.700 1154.310 1511.300 ;
      RECT 1156.270 0.700 1156.550 1511.300 ;
      RECT 1158.510 0.700 1158.790 1511.300 ;
      RECT 1160.750 0.700 1161.030 1511.300 ;
      RECT 1162.990 0.700 1163.270 1511.300 ;
      RECT 1165.230 0.700 1165.510 1511.300 ;
      RECT 1167.470 0.700 1167.750 1511.300 ;
      RECT 1169.710 0.700 1169.990 1511.300 ;
      RECT 1171.950 0.700 1172.230 1511.300 ;
      RECT 1174.190 0.700 1174.470 1511.300 ;
      RECT 1176.430 0.700 1176.710 1511.300 ;
      RECT 1178.670 0.700 1178.950 1511.300 ;
      RECT 1180.910 0.700 1181.190 1511.300 ;
      RECT 1183.150 0.700 1183.430 1511.300 ;
      RECT 1185.390 0.700 1185.670 1511.300 ;
      RECT 1187.630 0.700 1187.910 1511.300 ;
      RECT 1189.870 0.700 1190.150 1511.300 ;
      RECT 1192.110 0.700 1192.390 1511.300 ;
      RECT 1194.350 0.700 1194.630 1511.300 ;
      RECT 1196.590 0.700 1196.870 1511.300 ;
      RECT 1198.830 0.700 1199.110 1511.300 ;
      RECT 1201.070 0.700 1201.350 1511.300 ;
      RECT 1203.310 0.700 1203.590 1511.300 ;
      RECT 1205.550 0.700 1205.830 1511.300 ;
      RECT 1207.790 0.700 1208.070 1511.300 ;
      RECT 1210.030 0.700 1210.310 1511.300 ;
      RECT 1212.270 0.700 1212.550 1511.300 ;
      RECT 1214.510 0.700 1214.790 1511.300 ;
      RECT 1216.750 0.700 1217.030 1511.300 ;
      RECT 1218.990 0.700 1219.270 1511.300 ;
      RECT 1221.230 0.700 1221.510 1511.300 ;
      RECT 1223.470 0.700 1223.750 1511.300 ;
      RECT 1225.710 0.700 1225.990 1511.300 ;
      RECT 1227.950 0.700 1228.230 1511.300 ;
      RECT 1230.190 0.700 1230.470 1511.300 ;
      RECT 1232.430 0.700 1232.710 1511.300 ;
      RECT 1234.670 0.700 1234.950 1511.300 ;
      RECT 1236.910 0.700 1237.190 1511.300 ;
      RECT 1239.150 0.700 1239.430 1511.300 ;
      RECT 1241.390 0.700 1241.670 1511.300 ;
      RECT 1243.630 0.700 1243.910 1511.300 ;
      RECT 1245.870 0.700 1246.150 1511.300 ;
      RECT 1248.110 0.700 1248.390 1511.300 ;
      RECT 1250.350 0.700 1250.630 1511.300 ;
      RECT 1252.590 0.700 1252.870 1511.300 ;
      RECT 1254.830 0.700 1255.110 1511.300 ;
      RECT 1257.070 0.700 1257.350 1511.300 ;
      RECT 1259.310 0.700 1259.590 1511.300 ;
      RECT 1261.550 0.700 1261.830 1511.300 ;
      RECT 1263.790 0.700 1264.070 1511.300 ;
      RECT 1266.030 0.700 1266.310 1511.300 ;
      RECT 1268.270 0.700 1268.550 1511.300 ;
      RECT 1270.510 0.700 1270.790 1511.300 ;
      RECT 1272.750 0.700 1273.030 1511.300 ;
      RECT 1274.990 0.700 1275.270 1511.300 ;
      RECT 1277.230 0.700 1277.510 1511.300 ;
      RECT 1279.470 0.700 1279.750 1511.300 ;
      RECT 1281.710 0.700 1281.990 1511.300 ;
      RECT 1283.950 0.700 1284.230 1511.300 ;
      RECT 1286.190 0.700 1286.470 1511.300 ;
      RECT 1288.430 0.700 1288.710 1511.300 ;
      RECT 1290.670 0.700 1290.950 1511.300 ;
      RECT 1292.910 0.700 1293.190 1511.300 ;
      RECT 1295.150 0.700 1295.430 1511.300 ;
      RECT 1297.390 0.700 1297.670 1511.300 ;
      RECT 1299.630 0.700 1299.910 1511.300 ;
      RECT 1301.870 0.700 1302.150 1511.300 ;
      RECT 1304.110 0.700 1304.390 1511.300 ;
      RECT 1306.350 0.700 1306.630 1511.300 ;
      RECT 1308.590 0.700 1308.870 1511.300 ;
      RECT 1310.830 0.700 1311.110 1511.300 ;
      RECT 1313.070 0.700 1313.350 1511.300 ;
      RECT 1315.310 0.700 1315.590 1511.300 ;
      RECT 1317.550 0.700 1317.830 1511.300 ;
      RECT 1319.790 0.700 1320.070 1511.300 ;
      RECT 1322.030 0.700 1322.310 1511.300 ;
      RECT 1324.270 0.700 1324.550 1511.300 ;
      RECT 1326.510 0.700 1326.790 1511.300 ;
      RECT 1328.750 0.700 1329.030 1511.300 ;
      RECT 1330.990 0.700 1331.270 1511.300 ;
      RECT 1333.230 0.700 1333.510 1511.300 ;
      RECT 1335.470 0.700 1335.750 1511.300 ;
      RECT 1337.710 0.700 1337.990 1511.300 ;
      RECT 1339.950 0.700 1340.230 1511.300 ;
      RECT 1342.190 0.700 1342.470 1511.300 ;
      RECT 1344.430 0.700 1344.710 1511.300 ;
      RECT 1346.670 0.700 1346.950 1511.300 ;
      RECT 1348.910 0.700 1349.190 1511.300 ;
      RECT 1351.150 0.700 1351.430 1511.300 ;
      RECT 1353.390 0.700 1353.670 1511.300 ;
      RECT 1355.630 0.700 1355.910 1511.300 ;
      RECT 1357.870 0.700 1358.150 1511.300 ;
      RECT 1360.110 0.700 1360.390 1511.300 ;
      RECT 1362.350 0.700 1362.630 1511.300 ;
      RECT 1364.590 0.700 1364.870 1511.300 ;
      RECT 1366.830 0.700 1367.110 1511.300 ;
      RECT 1369.070 0.700 1369.350 1511.300 ;
      RECT 1371.310 0.700 1371.590 1511.300 ;
      RECT 1373.550 0.700 1373.830 1511.300 ;
      RECT 1375.790 0.700 1376.070 1511.300 ;
      RECT 1378.030 0.700 1378.310 1511.300 ;
      RECT 1380.270 0.700 1380.550 1511.300 ;
      RECT 1382.510 0.700 1382.790 1511.300 ;
      RECT 1384.750 0.700 1385.030 1511.300 ;
      RECT 1386.990 0.700 1387.270 1511.300 ;
      RECT 1389.230 0.700 1389.510 1511.300 ;
      RECT 1391.470 0.700 1391.750 1511.300 ;
      RECT 1393.710 0.700 1393.990 1511.300 ;
      RECT 1395.950 0.700 1396.230 1511.300 ;
      RECT 1398.190 0.700 1398.470 1511.300 ;
      RECT 1400.430 0.700 1400.710 1511.300 ;
      RECT 1402.670 0.700 1402.950 1511.300 ;
      RECT 1404.910 0.700 1405.190 1511.300 ;
      RECT 1407.150 0.700 1407.430 1511.300 ;
      RECT 1409.390 0.700 1409.670 1511.300 ;
      RECT 1411.630 0.700 1411.910 1511.300 ;
      RECT 1413.870 0.700 1414.150 1511.300 ;
      RECT 1416.110 0.700 1416.390 1511.300 ;
      RECT 1418.350 0.700 1418.630 1511.300 ;
      RECT 1420.590 0.700 1420.870 1511.300 ;
      RECT 1422.830 0.700 1423.110 1511.300 ;
      RECT 1425.070 0.700 1425.350 1511.300 ;
      RECT 1427.310 0.700 1427.590 1511.300 ;
      RECT 1429.550 0.700 1429.830 1511.300 ;
      RECT 1431.790 0.700 1432.070 1511.300 ;
      RECT 1434.030 0.700 1434.310 1511.300 ;
      RECT 1436.270 0.700 1436.550 1511.300 ;
      RECT 1438.510 0.700 1438.790 1511.300 ;
      RECT 1440.750 0.700 1441.030 1511.300 ;
      RECT 1442.990 0.700 1443.270 1511.300 ;
      RECT 1445.230 0.700 1445.510 1511.300 ;
      RECT 1447.470 0.700 1447.750 1511.300 ;
      RECT 1449.710 0.700 1449.990 1511.300 ;
      RECT 1451.950 0.700 1452.230 1511.300 ;
      RECT 1454.190 0.700 1454.470 1511.300 ;
      RECT 1456.430 0.700 1456.710 1511.300 ;
      RECT 1458.670 0.700 1458.950 1511.300 ;
      RECT 1460.910 0.700 1461.190 1511.300 ;
      RECT 1463.150 0.700 1463.430 1511.300 ;
      RECT 1465.390 0.700 1465.670 1511.300 ;
      RECT 1467.630 0.700 1467.910 1511.300 ;
      RECT 1469.870 0.700 1470.150 1511.300 ;
      RECT 1472.110 0.700 1472.390 1511.300 ;
      RECT 1474.350 0.700 1474.630 1511.300 ;
      RECT 1476.590 0.700 1476.870 1511.300 ;
      RECT 1478.830 0.700 1479.110 1511.300 ;
      RECT 1481.070 0.700 1481.350 1511.300 ;
      RECT 1483.310 0.700 1483.590 1511.300 ;
      RECT 1485.550 0.700 1485.830 1511.300 ;
      RECT 1487.790 0.700 1488.070 1511.300 ;
      RECT 1490.030 0.700 1490.310 1511.300 ;
      RECT 1492.270 0.700 1492.550 1511.300 ;
      RECT 1494.510 0.700 1494.790 1511.300 ;
      RECT 1496.750 0.700 1497.030 1511.300 ;
      RECT 1498.990 0.700 1499.270 1511.300 ;
      RECT 1501.230 0.700 1501.510 1511.300 ;
      RECT 1503.470 0.700 1503.750 1511.300 ;
      RECT 1505.710 0.700 1505.990 1511.300 ;
      RECT 1507.950 0.700 1508.230 1511.300 ;
      RECT 1510.190 0.700 1510.470 1511.300 ;
      RECT 1512.430 0.700 1512.710 1511.300 ;
      RECT 1514.670 0.700 1514.950 1511.300 ;
      RECT 1516.910 0.700 1517.190 1511.300 ;
      RECT 1519.150 0.700 1519.430 1511.300 ;
      RECT 1521.390 0.700 1521.670 1511.300 ;
      RECT 1523.630 0.700 1523.910 1511.300 ;
      RECT 1525.870 0.700 1526.150 1511.300 ;
      RECT 1528.110 0.700 1528.390 1511.300 ;
      RECT 1530.350 0.700 1530.630 1511.300 ;
      RECT 1532.590 0.700 1532.870 1511.300 ;
      RECT 1534.830 0.700 1535.110 1511.300 ;
      RECT 1537.070 0.700 1537.350 1511.300 ;
      RECT 1539.310 0.700 1539.590 1511.300 ;
      RECT 1541.550 0.700 1541.830 1511.300 ;
      RECT 1543.790 0.700 1544.070 1511.300 ;
      RECT 1546.030 0.700 1546.310 1511.300 ;
      RECT 1548.270 0.700 1548.550 1511.300 ;
      RECT 1550.510 0.700 1550.790 1511.300 ;
      RECT 1552.750 0.700 1553.030 1511.300 ;
      RECT 1554.990 0.700 1555.270 1511.300 ;
      RECT 1557.230 0.700 1557.510 1511.300 ;
      RECT 1559.470 0.700 1559.750 1511.300 ;
      RECT 1561.710 0.700 1561.990 1511.300 ;
      RECT 1563.950 0.700 1564.230 1511.300 ;
      RECT 1566.190 0.700 1566.470 1511.300 ;
      RECT 1568.430 0.700 1568.710 1511.300 ;
      RECT 1570.670 0.700 1570.950 1511.300 ;
      RECT 1572.910 0.700 1573.190 1511.300 ;
      RECT 1575.150 0.700 1575.430 1511.300 ;
      RECT 1577.390 0.700 1577.670 1511.300 ;
      RECT 1579.630 0.700 1579.910 1511.300 ;
      RECT 1581.870 0.700 1582.150 1511.300 ;
      RECT 1584.110 0.700 1584.390 1511.300 ;
      RECT 1586.350 0.700 1586.630 1511.300 ;
      RECT 1588.590 0.700 1588.870 1511.300 ;
      RECT 1590.830 0.700 1591.110 1511.300 ;
      RECT 1593.070 0.700 1593.350 1511.300 ;
      RECT 1595.310 0.700 1595.590 1511.300 ;
      RECT 1597.550 0.700 1597.830 1511.300 ;
      RECT 1599.790 0.700 1600.070 1511.300 ;
      RECT 1602.030 0.700 1602.310 1511.300 ;
      RECT 1604.270 0.700 1604.550 1511.300 ;
      RECT 1606.510 0.700 1606.790 1511.300 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 0.430 0.700 0.710 1511.300 ;
      RECT 2.670 0.700 2.950 1511.300 ;
      RECT 4.910 0.700 5.190 1511.300 ;
      RECT 7.150 0.700 7.430 1511.300 ;
      RECT 9.390 0.700 9.670 1511.300 ;
      RECT 11.630 0.700 11.910 1511.300 ;
      RECT 13.870 0.700 14.150 1511.300 ;
      RECT 16.110 0.700 16.390 1511.300 ;
      RECT 18.350 0.700 18.630 1511.300 ;
      RECT 20.590 0.700 20.870 1511.300 ;
      RECT 22.830 0.700 23.110 1511.300 ;
      RECT 25.070 0.700 25.350 1511.300 ;
      RECT 27.310 0.700 27.590 1511.300 ;
      RECT 29.550 0.700 29.830 1511.300 ;
      RECT 31.790 0.700 32.070 1511.300 ;
      RECT 34.030 0.700 34.310 1511.300 ;
      RECT 36.270 0.700 36.550 1511.300 ;
      RECT 38.510 0.700 38.790 1511.300 ;
      RECT 40.750 0.700 41.030 1511.300 ;
      RECT 42.990 0.700 43.270 1511.300 ;
      RECT 45.230 0.700 45.510 1511.300 ;
      RECT 47.470 0.700 47.750 1511.300 ;
      RECT 49.710 0.700 49.990 1511.300 ;
      RECT 51.950 0.700 52.230 1511.300 ;
      RECT 54.190 0.700 54.470 1511.300 ;
      RECT 56.430 0.700 56.710 1511.300 ;
      RECT 58.670 0.700 58.950 1511.300 ;
      RECT 60.910 0.700 61.190 1511.300 ;
      RECT 63.150 0.700 63.430 1511.300 ;
      RECT 65.390 0.700 65.670 1511.300 ;
      RECT 67.630 0.700 67.910 1511.300 ;
      RECT 69.870 0.700 70.150 1511.300 ;
      RECT 72.110 0.700 72.390 1511.300 ;
      RECT 74.350 0.700 74.630 1511.300 ;
      RECT 76.590 0.700 76.870 1511.300 ;
      RECT 78.830 0.700 79.110 1511.300 ;
      RECT 81.070 0.700 81.350 1511.300 ;
      RECT 83.310 0.700 83.590 1511.300 ;
      RECT 85.550 0.700 85.830 1511.300 ;
      RECT 87.790 0.700 88.070 1511.300 ;
      RECT 90.030 0.700 90.310 1511.300 ;
      RECT 92.270 0.700 92.550 1511.300 ;
      RECT 94.510 0.700 94.790 1511.300 ;
      RECT 96.750 0.700 97.030 1511.300 ;
      RECT 98.990 0.700 99.270 1511.300 ;
      RECT 101.230 0.700 101.510 1511.300 ;
      RECT 103.470 0.700 103.750 1511.300 ;
      RECT 105.710 0.700 105.990 1511.300 ;
      RECT 107.950 0.700 108.230 1511.300 ;
      RECT 110.190 0.700 110.470 1511.300 ;
      RECT 112.430 0.700 112.710 1511.300 ;
      RECT 114.670 0.700 114.950 1511.300 ;
      RECT 116.910 0.700 117.190 1511.300 ;
      RECT 119.150 0.700 119.430 1511.300 ;
      RECT 121.390 0.700 121.670 1511.300 ;
      RECT 123.630 0.700 123.910 1511.300 ;
      RECT 125.870 0.700 126.150 1511.300 ;
      RECT 128.110 0.700 128.390 1511.300 ;
      RECT 130.350 0.700 130.630 1511.300 ;
      RECT 132.590 0.700 132.870 1511.300 ;
      RECT 134.830 0.700 135.110 1511.300 ;
      RECT 137.070 0.700 137.350 1511.300 ;
      RECT 139.310 0.700 139.590 1511.300 ;
      RECT 141.550 0.700 141.830 1511.300 ;
      RECT 143.790 0.700 144.070 1511.300 ;
      RECT 146.030 0.700 146.310 1511.300 ;
      RECT 148.270 0.700 148.550 1511.300 ;
      RECT 150.510 0.700 150.790 1511.300 ;
      RECT 152.750 0.700 153.030 1511.300 ;
      RECT 154.990 0.700 155.270 1511.300 ;
      RECT 157.230 0.700 157.510 1511.300 ;
      RECT 159.470 0.700 159.750 1511.300 ;
      RECT 161.710 0.700 161.990 1511.300 ;
      RECT 163.950 0.700 164.230 1511.300 ;
      RECT 166.190 0.700 166.470 1511.300 ;
      RECT 168.430 0.700 168.710 1511.300 ;
      RECT 170.670 0.700 170.950 1511.300 ;
      RECT 172.910 0.700 173.190 1511.300 ;
      RECT 175.150 0.700 175.430 1511.300 ;
      RECT 177.390 0.700 177.670 1511.300 ;
      RECT 179.630 0.700 179.910 1511.300 ;
      RECT 181.870 0.700 182.150 1511.300 ;
      RECT 184.110 0.700 184.390 1511.300 ;
      RECT 186.350 0.700 186.630 1511.300 ;
      RECT 188.590 0.700 188.870 1511.300 ;
      RECT 190.830 0.700 191.110 1511.300 ;
      RECT 193.070 0.700 193.350 1511.300 ;
      RECT 195.310 0.700 195.590 1511.300 ;
      RECT 197.550 0.700 197.830 1511.300 ;
      RECT 199.790 0.700 200.070 1511.300 ;
      RECT 202.030 0.700 202.310 1511.300 ;
      RECT 204.270 0.700 204.550 1511.300 ;
      RECT 206.510 0.700 206.790 1511.300 ;
      RECT 208.750 0.700 209.030 1511.300 ;
      RECT 210.990 0.700 211.270 1511.300 ;
      RECT 213.230 0.700 213.510 1511.300 ;
      RECT 215.470 0.700 215.750 1511.300 ;
      RECT 217.710 0.700 217.990 1511.300 ;
      RECT 219.950 0.700 220.230 1511.300 ;
      RECT 222.190 0.700 222.470 1511.300 ;
      RECT 224.430 0.700 224.710 1511.300 ;
      RECT 226.670 0.700 226.950 1511.300 ;
      RECT 228.910 0.700 229.190 1511.300 ;
      RECT 231.150 0.700 231.430 1511.300 ;
      RECT 233.390 0.700 233.670 1511.300 ;
      RECT 235.630 0.700 235.910 1511.300 ;
      RECT 237.870 0.700 238.150 1511.300 ;
      RECT 240.110 0.700 240.390 1511.300 ;
      RECT 242.350 0.700 242.630 1511.300 ;
      RECT 244.590 0.700 244.870 1511.300 ;
      RECT 246.830 0.700 247.110 1511.300 ;
      RECT 249.070 0.700 249.350 1511.300 ;
      RECT 251.310 0.700 251.590 1511.300 ;
      RECT 253.550 0.700 253.830 1511.300 ;
      RECT 255.790 0.700 256.070 1511.300 ;
      RECT 258.030 0.700 258.310 1511.300 ;
      RECT 260.270 0.700 260.550 1511.300 ;
      RECT 262.510 0.700 262.790 1511.300 ;
      RECT 264.750 0.700 265.030 1511.300 ;
      RECT 266.990 0.700 267.270 1511.300 ;
      RECT 269.230 0.700 269.510 1511.300 ;
      RECT 271.470 0.700 271.750 1511.300 ;
      RECT 273.710 0.700 273.990 1511.300 ;
      RECT 275.950 0.700 276.230 1511.300 ;
      RECT 278.190 0.700 278.470 1511.300 ;
      RECT 280.430 0.700 280.710 1511.300 ;
      RECT 282.670 0.700 282.950 1511.300 ;
      RECT 284.910 0.700 285.190 1511.300 ;
      RECT 287.150 0.700 287.430 1511.300 ;
      RECT 289.390 0.700 289.670 1511.300 ;
      RECT 291.630 0.700 291.910 1511.300 ;
      RECT 293.870 0.700 294.150 1511.300 ;
      RECT 296.110 0.700 296.390 1511.300 ;
      RECT 298.350 0.700 298.630 1511.300 ;
      RECT 300.590 0.700 300.870 1511.300 ;
      RECT 302.830 0.700 303.110 1511.300 ;
      RECT 305.070 0.700 305.350 1511.300 ;
      RECT 307.310 0.700 307.590 1511.300 ;
      RECT 309.550 0.700 309.830 1511.300 ;
      RECT 311.790 0.700 312.070 1511.300 ;
      RECT 314.030 0.700 314.310 1511.300 ;
      RECT 316.270 0.700 316.550 1511.300 ;
      RECT 318.510 0.700 318.790 1511.300 ;
      RECT 320.750 0.700 321.030 1511.300 ;
      RECT 322.990 0.700 323.270 1511.300 ;
      RECT 325.230 0.700 325.510 1511.300 ;
      RECT 327.470 0.700 327.750 1511.300 ;
      RECT 329.710 0.700 329.990 1511.300 ;
      RECT 331.950 0.700 332.230 1511.300 ;
      RECT 334.190 0.700 334.470 1511.300 ;
      RECT 336.430 0.700 336.710 1511.300 ;
      RECT 338.670 0.700 338.950 1511.300 ;
      RECT 340.910 0.700 341.190 1511.300 ;
      RECT 343.150 0.700 343.430 1511.300 ;
      RECT 345.390 0.700 345.670 1511.300 ;
      RECT 347.630 0.700 347.910 1511.300 ;
      RECT 349.870 0.700 350.150 1511.300 ;
      RECT 352.110 0.700 352.390 1511.300 ;
      RECT 354.350 0.700 354.630 1511.300 ;
      RECT 356.590 0.700 356.870 1511.300 ;
      RECT 358.830 0.700 359.110 1511.300 ;
      RECT 361.070 0.700 361.350 1511.300 ;
      RECT 363.310 0.700 363.590 1511.300 ;
      RECT 365.550 0.700 365.830 1511.300 ;
      RECT 367.790 0.700 368.070 1511.300 ;
      RECT 370.030 0.700 370.310 1511.300 ;
      RECT 372.270 0.700 372.550 1511.300 ;
      RECT 374.510 0.700 374.790 1511.300 ;
      RECT 376.750 0.700 377.030 1511.300 ;
      RECT 378.990 0.700 379.270 1511.300 ;
      RECT 381.230 0.700 381.510 1511.300 ;
      RECT 383.470 0.700 383.750 1511.300 ;
      RECT 385.710 0.700 385.990 1511.300 ;
      RECT 387.950 0.700 388.230 1511.300 ;
      RECT 390.190 0.700 390.470 1511.300 ;
      RECT 392.430 0.700 392.710 1511.300 ;
      RECT 394.670 0.700 394.950 1511.300 ;
      RECT 396.910 0.700 397.190 1511.300 ;
      RECT 399.150 0.700 399.430 1511.300 ;
      RECT 401.390 0.700 401.670 1511.300 ;
      RECT 403.630 0.700 403.910 1511.300 ;
      RECT 405.870 0.700 406.150 1511.300 ;
      RECT 408.110 0.700 408.390 1511.300 ;
      RECT 410.350 0.700 410.630 1511.300 ;
      RECT 412.590 0.700 412.870 1511.300 ;
      RECT 414.830 0.700 415.110 1511.300 ;
      RECT 417.070 0.700 417.350 1511.300 ;
      RECT 419.310 0.700 419.590 1511.300 ;
      RECT 421.550 0.700 421.830 1511.300 ;
      RECT 423.790 0.700 424.070 1511.300 ;
      RECT 426.030 0.700 426.310 1511.300 ;
      RECT 428.270 0.700 428.550 1511.300 ;
      RECT 430.510 0.700 430.790 1511.300 ;
      RECT 432.750 0.700 433.030 1511.300 ;
      RECT 434.990 0.700 435.270 1511.300 ;
      RECT 437.230 0.700 437.510 1511.300 ;
      RECT 439.470 0.700 439.750 1511.300 ;
      RECT 441.710 0.700 441.990 1511.300 ;
      RECT 443.950 0.700 444.230 1511.300 ;
      RECT 446.190 0.700 446.470 1511.300 ;
      RECT 448.430 0.700 448.710 1511.300 ;
      RECT 450.670 0.700 450.950 1511.300 ;
      RECT 452.910 0.700 453.190 1511.300 ;
      RECT 455.150 0.700 455.430 1511.300 ;
      RECT 457.390 0.700 457.670 1511.300 ;
      RECT 459.630 0.700 459.910 1511.300 ;
      RECT 461.870 0.700 462.150 1511.300 ;
      RECT 464.110 0.700 464.390 1511.300 ;
      RECT 466.350 0.700 466.630 1511.300 ;
      RECT 468.590 0.700 468.870 1511.300 ;
      RECT 470.830 0.700 471.110 1511.300 ;
      RECT 473.070 0.700 473.350 1511.300 ;
      RECT 475.310 0.700 475.590 1511.300 ;
      RECT 477.550 0.700 477.830 1511.300 ;
      RECT 479.790 0.700 480.070 1511.300 ;
      RECT 482.030 0.700 482.310 1511.300 ;
      RECT 484.270 0.700 484.550 1511.300 ;
      RECT 486.510 0.700 486.790 1511.300 ;
      RECT 488.750 0.700 489.030 1511.300 ;
      RECT 490.990 0.700 491.270 1511.300 ;
      RECT 493.230 0.700 493.510 1511.300 ;
      RECT 495.470 0.700 495.750 1511.300 ;
      RECT 497.710 0.700 497.990 1511.300 ;
      RECT 499.950 0.700 500.230 1511.300 ;
      RECT 502.190 0.700 502.470 1511.300 ;
      RECT 504.430 0.700 504.710 1511.300 ;
      RECT 506.670 0.700 506.950 1511.300 ;
      RECT 508.910 0.700 509.190 1511.300 ;
      RECT 511.150 0.700 511.430 1511.300 ;
      RECT 513.390 0.700 513.670 1511.300 ;
      RECT 515.630 0.700 515.910 1511.300 ;
      RECT 517.870 0.700 518.150 1511.300 ;
      RECT 520.110 0.700 520.390 1511.300 ;
      RECT 522.350 0.700 522.630 1511.300 ;
      RECT 524.590 0.700 524.870 1511.300 ;
      RECT 526.830 0.700 527.110 1511.300 ;
      RECT 529.070 0.700 529.350 1511.300 ;
      RECT 531.310 0.700 531.590 1511.300 ;
      RECT 533.550 0.700 533.830 1511.300 ;
      RECT 535.790 0.700 536.070 1511.300 ;
      RECT 538.030 0.700 538.310 1511.300 ;
      RECT 540.270 0.700 540.550 1511.300 ;
      RECT 542.510 0.700 542.790 1511.300 ;
      RECT 544.750 0.700 545.030 1511.300 ;
      RECT 546.990 0.700 547.270 1511.300 ;
      RECT 549.230 0.700 549.510 1511.300 ;
      RECT 551.470 0.700 551.750 1511.300 ;
      RECT 553.710 0.700 553.990 1511.300 ;
      RECT 555.950 0.700 556.230 1511.300 ;
      RECT 558.190 0.700 558.470 1511.300 ;
      RECT 560.430 0.700 560.710 1511.300 ;
      RECT 562.670 0.700 562.950 1511.300 ;
      RECT 564.910 0.700 565.190 1511.300 ;
      RECT 567.150 0.700 567.430 1511.300 ;
      RECT 569.390 0.700 569.670 1511.300 ;
      RECT 571.630 0.700 571.910 1511.300 ;
      RECT 573.870 0.700 574.150 1511.300 ;
      RECT 576.110 0.700 576.390 1511.300 ;
      RECT 578.350 0.700 578.630 1511.300 ;
      RECT 580.590 0.700 580.870 1511.300 ;
      RECT 582.830 0.700 583.110 1511.300 ;
      RECT 585.070 0.700 585.350 1511.300 ;
      RECT 587.310 0.700 587.590 1511.300 ;
      RECT 589.550 0.700 589.830 1511.300 ;
      RECT 591.790 0.700 592.070 1511.300 ;
      RECT 594.030 0.700 594.310 1511.300 ;
      RECT 596.270 0.700 596.550 1511.300 ;
      RECT 598.510 0.700 598.790 1511.300 ;
      RECT 600.750 0.700 601.030 1511.300 ;
      RECT 602.990 0.700 603.270 1511.300 ;
      RECT 605.230 0.700 605.510 1511.300 ;
      RECT 607.470 0.700 607.750 1511.300 ;
      RECT 609.710 0.700 609.990 1511.300 ;
      RECT 611.950 0.700 612.230 1511.300 ;
      RECT 614.190 0.700 614.470 1511.300 ;
      RECT 616.430 0.700 616.710 1511.300 ;
      RECT 618.670 0.700 618.950 1511.300 ;
      RECT 620.910 0.700 621.190 1511.300 ;
      RECT 623.150 0.700 623.430 1511.300 ;
      RECT 625.390 0.700 625.670 1511.300 ;
      RECT 627.630 0.700 627.910 1511.300 ;
      RECT 629.870 0.700 630.150 1511.300 ;
      RECT 632.110 0.700 632.390 1511.300 ;
      RECT 634.350 0.700 634.630 1511.300 ;
      RECT 636.590 0.700 636.870 1511.300 ;
      RECT 638.830 0.700 639.110 1511.300 ;
      RECT 641.070 0.700 641.350 1511.300 ;
      RECT 643.310 0.700 643.590 1511.300 ;
      RECT 645.550 0.700 645.830 1511.300 ;
      RECT 647.790 0.700 648.070 1511.300 ;
      RECT 650.030 0.700 650.310 1511.300 ;
      RECT 652.270 0.700 652.550 1511.300 ;
      RECT 654.510 0.700 654.790 1511.300 ;
      RECT 656.750 0.700 657.030 1511.300 ;
      RECT 658.990 0.700 659.270 1511.300 ;
      RECT 661.230 0.700 661.510 1511.300 ;
      RECT 663.470 0.700 663.750 1511.300 ;
      RECT 665.710 0.700 665.990 1511.300 ;
      RECT 667.950 0.700 668.230 1511.300 ;
      RECT 670.190 0.700 670.470 1511.300 ;
      RECT 672.430 0.700 672.710 1511.300 ;
      RECT 674.670 0.700 674.950 1511.300 ;
      RECT 676.910 0.700 677.190 1511.300 ;
      RECT 679.150 0.700 679.430 1511.300 ;
      RECT 681.390 0.700 681.670 1511.300 ;
      RECT 683.630 0.700 683.910 1511.300 ;
      RECT 685.870 0.700 686.150 1511.300 ;
      RECT 688.110 0.700 688.390 1511.300 ;
      RECT 690.350 0.700 690.630 1511.300 ;
      RECT 692.590 0.700 692.870 1511.300 ;
      RECT 694.830 0.700 695.110 1511.300 ;
      RECT 697.070 0.700 697.350 1511.300 ;
      RECT 699.310 0.700 699.590 1511.300 ;
      RECT 701.550 0.700 701.830 1511.300 ;
      RECT 703.790 0.700 704.070 1511.300 ;
      RECT 706.030 0.700 706.310 1511.300 ;
      RECT 708.270 0.700 708.550 1511.300 ;
      RECT 710.510 0.700 710.790 1511.300 ;
      RECT 712.750 0.700 713.030 1511.300 ;
      RECT 714.990 0.700 715.270 1511.300 ;
      RECT 717.230 0.700 717.510 1511.300 ;
      RECT 719.470 0.700 719.750 1511.300 ;
      RECT 721.710 0.700 721.990 1511.300 ;
      RECT 723.950 0.700 724.230 1511.300 ;
      RECT 726.190 0.700 726.470 1511.300 ;
      RECT 728.430 0.700 728.710 1511.300 ;
      RECT 730.670 0.700 730.950 1511.300 ;
      RECT 732.910 0.700 733.190 1511.300 ;
      RECT 735.150 0.700 735.430 1511.300 ;
      RECT 737.390 0.700 737.670 1511.300 ;
      RECT 739.630 0.700 739.910 1511.300 ;
      RECT 741.870 0.700 742.150 1511.300 ;
      RECT 744.110 0.700 744.390 1511.300 ;
      RECT 746.350 0.700 746.630 1511.300 ;
      RECT 748.590 0.700 748.870 1511.300 ;
      RECT 750.830 0.700 751.110 1511.300 ;
      RECT 753.070 0.700 753.350 1511.300 ;
      RECT 755.310 0.700 755.590 1511.300 ;
      RECT 757.550 0.700 757.830 1511.300 ;
      RECT 759.790 0.700 760.070 1511.300 ;
      RECT 762.030 0.700 762.310 1511.300 ;
      RECT 764.270 0.700 764.550 1511.300 ;
      RECT 766.510 0.700 766.790 1511.300 ;
      RECT 768.750 0.700 769.030 1511.300 ;
      RECT 770.990 0.700 771.270 1511.300 ;
      RECT 773.230 0.700 773.510 1511.300 ;
      RECT 775.470 0.700 775.750 1511.300 ;
      RECT 777.710 0.700 777.990 1511.300 ;
      RECT 779.950 0.700 780.230 1511.300 ;
      RECT 782.190 0.700 782.470 1511.300 ;
      RECT 784.430 0.700 784.710 1511.300 ;
      RECT 786.670 0.700 786.950 1511.300 ;
      RECT 788.910 0.700 789.190 1511.300 ;
      RECT 791.150 0.700 791.430 1511.300 ;
      RECT 793.390 0.700 793.670 1511.300 ;
      RECT 795.630 0.700 795.910 1511.300 ;
      RECT 797.870 0.700 798.150 1511.300 ;
      RECT 800.110 0.700 800.390 1511.300 ;
      RECT 802.350 0.700 802.630 1511.300 ;
      RECT 804.590 0.700 804.870 1511.300 ;
      RECT 806.830 0.700 807.110 1511.300 ;
      RECT 809.070 0.700 809.350 1511.300 ;
      RECT 811.310 0.700 811.590 1511.300 ;
      RECT 813.550 0.700 813.830 1511.300 ;
      RECT 815.790 0.700 816.070 1511.300 ;
      RECT 818.030 0.700 818.310 1511.300 ;
      RECT 820.270 0.700 820.550 1511.300 ;
      RECT 822.510 0.700 822.790 1511.300 ;
      RECT 824.750 0.700 825.030 1511.300 ;
      RECT 826.990 0.700 827.270 1511.300 ;
      RECT 829.230 0.700 829.510 1511.300 ;
      RECT 831.470 0.700 831.750 1511.300 ;
      RECT 833.710 0.700 833.990 1511.300 ;
      RECT 835.950 0.700 836.230 1511.300 ;
      RECT 838.190 0.700 838.470 1511.300 ;
      RECT 840.430 0.700 840.710 1511.300 ;
      RECT 842.670 0.700 842.950 1511.300 ;
      RECT 844.910 0.700 845.190 1511.300 ;
      RECT 847.150 0.700 847.430 1511.300 ;
      RECT 849.390 0.700 849.670 1511.300 ;
      RECT 851.630 0.700 851.910 1511.300 ;
      RECT 853.870 0.700 854.150 1511.300 ;
      RECT 856.110 0.700 856.390 1511.300 ;
      RECT 858.350 0.700 858.630 1511.300 ;
      RECT 860.590 0.700 860.870 1511.300 ;
      RECT 862.830 0.700 863.110 1511.300 ;
      RECT 865.070 0.700 865.350 1511.300 ;
      RECT 867.310 0.700 867.590 1511.300 ;
      RECT 869.550 0.700 869.830 1511.300 ;
      RECT 871.790 0.700 872.070 1511.300 ;
      RECT 874.030 0.700 874.310 1511.300 ;
      RECT 876.270 0.700 876.550 1511.300 ;
      RECT 878.510 0.700 878.790 1511.300 ;
      RECT 880.750 0.700 881.030 1511.300 ;
      RECT 882.990 0.700 883.270 1511.300 ;
      RECT 885.230 0.700 885.510 1511.300 ;
      RECT 887.470 0.700 887.750 1511.300 ;
      RECT 889.710 0.700 889.990 1511.300 ;
      RECT 891.950 0.700 892.230 1511.300 ;
      RECT 894.190 0.700 894.470 1511.300 ;
      RECT 896.430 0.700 896.710 1511.300 ;
      RECT 898.670 0.700 898.950 1511.300 ;
      RECT 900.910 0.700 901.190 1511.300 ;
      RECT 903.150 0.700 903.430 1511.300 ;
      RECT 905.390 0.700 905.670 1511.300 ;
      RECT 907.630 0.700 907.910 1511.300 ;
      RECT 909.870 0.700 910.150 1511.300 ;
      RECT 912.110 0.700 912.390 1511.300 ;
      RECT 914.350 0.700 914.630 1511.300 ;
      RECT 916.590 0.700 916.870 1511.300 ;
      RECT 918.830 0.700 919.110 1511.300 ;
      RECT 921.070 0.700 921.350 1511.300 ;
      RECT 923.310 0.700 923.590 1511.300 ;
      RECT 925.550 0.700 925.830 1511.300 ;
      RECT 927.790 0.700 928.070 1511.300 ;
      RECT 930.030 0.700 930.310 1511.300 ;
      RECT 932.270 0.700 932.550 1511.300 ;
      RECT 934.510 0.700 934.790 1511.300 ;
      RECT 936.750 0.700 937.030 1511.300 ;
      RECT 938.990 0.700 939.270 1511.300 ;
      RECT 941.230 0.700 941.510 1511.300 ;
      RECT 943.470 0.700 943.750 1511.300 ;
      RECT 945.710 0.700 945.990 1511.300 ;
      RECT 947.950 0.700 948.230 1511.300 ;
      RECT 950.190 0.700 950.470 1511.300 ;
      RECT 952.430 0.700 952.710 1511.300 ;
      RECT 954.670 0.700 954.950 1511.300 ;
      RECT 956.910 0.700 957.190 1511.300 ;
      RECT 959.150 0.700 959.430 1511.300 ;
      RECT 961.390 0.700 961.670 1511.300 ;
      RECT 963.630 0.700 963.910 1511.300 ;
      RECT 965.870 0.700 966.150 1511.300 ;
      RECT 968.110 0.700 968.390 1511.300 ;
      RECT 970.350 0.700 970.630 1511.300 ;
      RECT 972.590 0.700 972.870 1511.300 ;
      RECT 974.830 0.700 975.110 1511.300 ;
      RECT 977.070 0.700 977.350 1511.300 ;
      RECT 979.310 0.700 979.590 1511.300 ;
      RECT 981.550 0.700 981.830 1511.300 ;
      RECT 983.790 0.700 984.070 1511.300 ;
      RECT 986.030 0.700 986.310 1511.300 ;
      RECT 988.270 0.700 988.550 1511.300 ;
      RECT 990.510 0.700 990.790 1511.300 ;
      RECT 992.750 0.700 993.030 1511.300 ;
      RECT 994.990 0.700 995.270 1511.300 ;
      RECT 997.230 0.700 997.510 1511.300 ;
      RECT 999.470 0.700 999.750 1511.300 ;
      RECT 1001.710 0.700 1001.990 1511.300 ;
      RECT 1003.950 0.700 1004.230 1511.300 ;
      RECT 1006.190 0.700 1006.470 1511.300 ;
      RECT 1008.430 0.700 1008.710 1511.300 ;
      RECT 1010.670 0.700 1010.950 1511.300 ;
      RECT 1012.910 0.700 1013.190 1511.300 ;
      RECT 1015.150 0.700 1015.430 1511.300 ;
      RECT 1017.390 0.700 1017.670 1511.300 ;
      RECT 1019.630 0.700 1019.910 1511.300 ;
      RECT 1021.870 0.700 1022.150 1511.300 ;
      RECT 1024.110 0.700 1024.390 1511.300 ;
      RECT 1026.350 0.700 1026.630 1511.300 ;
      RECT 1028.590 0.700 1028.870 1511.300 ;
      RECT 1030.830 0.700 1031.110 1511.300 ;
      RECT 1033.070 0.700 1033.350 1511.300 ;
      RECT 1035.310 0.700 1035.590 1511.300 ;
      RECT 1037.550 0.700 1037.830 1511.300 ;
      RECT 1039.790 0.700 1040.070 1511.300 ;
      RECT 1042.030 0.700 1042.310 1511.300 ;
      RECT 1044.270 0.700 1044.550 1511.300 ;
      RECT 1046.510 0.700 1046.790 1511.300 ;
      RECT 1048.750 0.700 1049.030 1511.300 ;
      RECT 1050.990 0.700 1051.270 1511.300 ;
      RECT 1053.230 0.700 1053.510 1511.300 ;
      RECT 1055.470 0.700 1055.750 1511.300 ;
      RECT 1057.710 0.700 1057.990 1511.300 ;
      RECT 1059.950 0.700 1060.230 1511.300 ;
      RECT 1062.190 0.700 1062.470 1511.300 ;
      RECT 1064.430 0.700 1064.710 1511.300 ;
      RECT 1066.670 0.700 1066.950 1511.300 ;
      RECT 1068.910 0.700 1069.190 1511.300 ;
      RECT 1071.150 0.700 1071.430 1511.300 ;
      RECT 1073.390 0.700 1073.670 1511.300 ;
      RECT 1075.630 0.700 1075.910 1511.300 ;
      RECT 1077.870 0.700 1078.150 1511.300 ;
      RECT 1080.110 0.700 1080.390 1511.300 ;
      RECT 1082.350 0.700 1082.630 1511.300 ;
      RECT 1084.590 0.700 1084.870 1511.300 ;
      RECT 1086.830 0.700 1087.110 1511.300 ;
      RECT 1089.070 0.700 1089.350 1511.300 ;
      RECT 1091.310 0.700 1091.590 1511.300 ;
      RECT 1093.550 0.700 1093.830 1511.300 ;
      RECT 1095.790 0.700 1096.070 1511.300 ;
      RECT 1098.030 0.700 1098.310 1511.300 ;
      RECT 1100.270 0.700 1100.550 1511.300 ;
      RECT 1102.510 0.700 1102.790 1511.300 ;
      RECT 1104.750 0.700 1105.030 1511.300 ;
      RECT 1106.990 0.700 1107.270 1511.300 ;
      RECT 1109.230 0.700 1109.510 1511.300 ;
      RECT 1111.470 0.700 1111.750 1511.300 ;
      RECT 1113.710 0.700 1113.990 1511.300 ;
      RECT 1115.950 0.700 1116.230 1511.300 ;
      RECT 1118.190 0.700 1118.470 1511.300 ;
      RECT 1120.430 0.700 1120.710 1511.300 ;
      RECT 1122.670 0.700 1122.950 1511.300 ;
      RECT 1124.910 0.700 1125.190 1511.300 ;
      RECT 1127.150 0.700 1127.430 1511.300 ;
      RECT 1129.390 0.700 1129.670 1511.300 ;
      RECT 1131.630 0.700 1131.910 1511.300 ;
      RECT 1133.870 0.700 1134.150 1511.300 ;
      RECT 1136.110 0.700 1136.390 1511.300 ;
      RECT 1138.350 0.700 1138.630 1511.300 ;
      RECT 1140.590 0.700 1140.870 1511.300 ;
      RECT 1142.830 0.700 1143.110 1511.300 ;
      RECT 1145.070 0.700 1145.350 1511.300 ;
      RECT 1147.310 0.700 1147.590 1511.300 ;
      RECT 1149.550 0.700 1149.830 1511.300 ;
      RECT 1151.790 0.700 1152.070 1511.300 ;
      RECT 1154.030 0.700 1154.310 1511.300 ;
      RECT 1156.270 0.700 1156.550 1511.300 ;
      RECT 1158.510 0.700 1158.790 1511.300 ;
      RECT 1160.750 0.700 1161.030 1511.300 ;
      RECT 1162.990 0.700 1163.270 1511.300 ;
      RECT 1165.230 0.700 1165.510 1511.300 ;
      RECT 1167.470 0.700 1167.750 1511.300 ;
      RECT 1169.710 0.700 1169.990 1511.300 ;
      RECT 1171.950 0.700 1172.230 1511.300 ;
      RECT 1174.190 0.700 1174.470 1511.300 ;
      RECT 1176.430 0.700 1176.710 1511.300 ;
      RECT 1178.670 0.700 1178.950 1511.300 ;
      RECT 1180.910 0.700 1181.190 1511.300 ;
      RECT 1183.150 0.700 1183.430 1511.300 ;
      RECT 1185.390 0.700 1185.670 1511.300 ;
      RECT 1187.630 0.700 1187.910 1511.300 ;
      RECT 1189.870 0.700 1190.150 1511.300 ;
      RECT 1192.110 0.700 1192.390 1511.300 ;
      RECT 1194.350 0.700 1194.630 1511.300 ;
      RECT 1196.590 0.700 1196.870 1511.300 ;
      RECT 1198.830 0.700 1199.110 1511.300 ;
      RECT 1201.070 0.700 1201.350 1511.300 ;
      RECT 1203.310 0.700 1203.590 1511.300 ;
      RECT 1205.550 0.700 1205.830 1511.300 ;
      RECT 1207.790 0.700 1208.070 1511.300 ;
      RECT 1210.030 0.700 1210.310 1511.300 ;
      RECT 1212.270 0.700 1212.550 1511.300 ;
      RECT 1214.510 0.700 1214.790 1511.300 ;
      RECT 1216.750 0.700 1217.030 1511.300 ;
      RECT 1218.990 0.700 1219.270 1511.300 ;
      RECT 1221.230 0.700 1221.510 1511.300 ;
      RECT 1223.470 0.700 1223.750 1511.300 ;
      RECT 1225.710 0.700 1225.990 1511.300 ;
      RECT 1227.950 0.700 1228.230 1511.300 ;
      RECT 1230.190 0.700 1230.470 1511.300 ;
      RECT 1232.430 0.700 1232.710 1511.300 ;
      RECT 1234.670 0.700 1234.950 1511.300 ;
      RECT 1236.910 0.700 1237.190 1511.300 ;
      RECT 1239.150 0.700 1239.430 1511.300 ;
      RECT 1241.390 0.700 1241.670 1511.300 ;
      RECT 1243.630 0.700 1243.910 1511.300 ;
      RECT 1245.870 0.700 1246.150 1511.300 ;
      RECT 1248.110 0.700 1248.390 1511.300 ;
      RECT 1250.350 0.700 1250.630 1511.300 ;
      RECT 1252.590 0.700 1252.870 1511.300 ;
      RECT 1254.830 0.700 1255.110 1511.300 ;
      RECT 1257.070 0.700 1257.350 1511.300 ;
      RECT 1259.310 0.700 1259.590 1511.300 ;
      RECT 1261.550 0.700 1261.830 1511.300 ;
      RECT 1263.790 0.700 1264.070 1511.300 ;
      RECT 1266.030 0.700 1266.310 1511.300 ;
      RECT 1268.270 0.700 1268.550 1511.300 ;
      RECT 1270.510 0.700 1270.790 1511.300 ;
      RECT 1272.750 0.700 1273.030 1511.300 ;
      RECT 1274.990 0.700 1275.270 1511.300 ;
      RECT 1277.230 0.700 1277.510 1511.300 ;
      RECT 1279.470 0.700 1279.750 1511.300 ;
      RECT 1281.710 0.700 1281.990 1511.300 ;
      RECT 1283.950 0.700 1284.230 1511.300 ;
      RECT 1286.190 0.700 1286.470 1511.300 ;
      RECT 1288.430 0.700 1288.710 1511.300 ;
      RECT 1290.670 0.700 1290.950 1511.300 ;
      RECT 1292.910 0.700 1293.190 1511.300 ;
      RECT 1295.150 0.700 1295.430 1511.300 ;
      RECT 1297.390 0.700 1297.670 1511.300 ;
      RECT 1299.630 0.700 1299.910 1511.300 ;
      RECT 1301.870 0.700 1302.150 1511.300 ;
      RECT 1304.110 0.700 1304.390 1511.300 ;
      RECT 1306.350 0.700 1306.630 1511.300 ;
      RECT 1308.590 0.700 1308.870 1511.300 ;
      RECT 1310.830 0.700 1311.110 1511.300 ;
      RECT 1313.070 0.700 1313.350 1511.300 ;
      RECT 1315.310 0.700 1315.590 1511.300 ;
      RECT 1317.550 0.700 1317.830 1511.300 ;
      RECT 1319.790 0.700 1320.070 1511.300 ;
      RECT 1322.030 0.700 1322.310 1511.300 ;
      RECT 1324.270 0.700 1324.550 1511.300 ;
      RECT 1326.510 0.700 1326.790 1511.300 ;
      RECT 1328.750 0.700 1329.030 1511.300 ;
      RECT 1330.990 0.700 1331.270 1511.300 ;
      RECT 1333.230 0.700 1333.510 1511.300 ;
      RECT 1335.470 0.700 1335.750 1511.300 ;
      RECT 1337.710 0.700 1337.990 1511.300 ;
      RECT 1339.950 0.700 1340.230 1511.300 ;
      RECT 1342.190 0.700 1342.470 1511.300 ;
      RECT 1344.430 0.700 1344.710 1511.300 ;
      RECT 1346.670 0.700 1346.950 1511.300 ;
      RECT 1348.910 0.700 1349.190 1511.300 ;
      RECT 1351.150 0.700 1351.430 1511.300 ;
      RECT 1353.390 0.700 1353.670 1511.300 ;
      RECT 1355.630 0.700 1355.910 1511.300 ;
      RECT 1357.870 0.700 1358.150 1511.300 ;
      RECT 1360.110 0.700 1360.390 1511.300 ;
      RECT 1362.350 0.700 1362.630 1511.300 ;
      RECT 1364.590 0.700 1364.870 1511.300 ;
      RECT 1366.830 0.700 1367.110 1511.300 ;
      RECT 1369.070 0.700 1369.350 1511.300 ;
      RECT 1371.310 0.700 1371.590 1511.300 ;
      RECT 1373.550 0.700 1373.830 1511.300 ;
      RECT 1375.790 0.700 1376.070 1511.300 ;
      RECT 1378.030 0.700 1378.310 1511.300 ;
      RECT 1380.270 0.700 1380.550 1511.300 ;
      RECT 1382.510 0.700 1382.790 1511.300 ;
      RECT 1384.750 0.700 1385.030 1511.300 ;
      RECT 1386.990 0.700 1387.270 1511.300 ;
      RECT 1389.230 0.700 1389.510 1511.300 ;
      RECT 1391.470 0.700 1391.750 1511.300 ;
      RECT 1393.710 0.700 1393.990 1511.300 ;
      RECT 1395.950 0.700 1396.230 1511.300 ;
      RECT 1398.190 0.700 1398.470 1511.300 ;
      RECT 1400.430 0.700 1400.710 1511.300 ;
      RECT 1402.670 0.700 1402.950 1511.300 ;
      RECT 1404.910 0.700 1405.190 1511.300 ;
      RECT 1407.150 0.700 1407.430 1511.300 ;
      RECT 1409.390 0.700 1409.670 1511.300 ;
      RECT 1411.630 0.700 1411.910 1511.300 ;
      RECT 1413.870 0.700 1414.150 1511.300 ;
      RECT 1416.110 0.700 1416.390 1511.300 ;
      RECT 1418.350 0.700 1418.630 1511.300 ;
      RECT 1420.590 0.700 1420.870 1511.300 ;
      RECT 1422.830 0.700 1423.110 1511.300 ;
      RECT 1425.070 0.700 1425.350 1511.300 ;
      RECT 1427.310 0.700 1427.590 1511.300 ;
      RECT 1429.550 0.700 1429.830 1511.300 ;
      RECT 1431.790 0.700 1432.070 1511.300 ;
      RECT 1434.030 0.700 1434.310 1511.300 ;
      RECT 1436.270 0.700 1436.550 1511.300 ;
      RECT 1438.510 0.700 1438.790 1511.300 ;
      RECT 1440.750 0.700 1441.030 1511.300 ;
      RECT 1442.990 0.700 1443.270 1511.300 ;
      RECT 1445.230 0.700 1445.510 1511.300 ;
      RECT 1447.470 0.700 1447.750 1511.300 ;
      RECT 1449.710 0.700 1449.990 1511.300 ;
      RECT 1451.950 0.700 1452.230 1511.300 ;
      RECT 1454.190 0.700 1454.470 1511.300 ;
      RECT 1456.430 0.700 1456.710 1511.300 ;
      RECT 1458.670 0.700 1458.950 1511.300 ;
      RECT 1460.910 0.700 1461.190 1511.300 ;
      RECT 1463.150 0.700 1463.430 1511.300 ;
      RECT 1465.390 0.700 1465.670 1511.300 ;
      RECT 1467.630 0.700 1467.910 1511.300 ;
      RECT 1469.870 0.700 1470.150 1511.300 ;
      RECT 1472.110 0.700 1472.390 1511.300 ;
      RECT 1474.350 0.700 1474.630 1511.300 ;
      RECT 1476.590 0.700 1476.870 1511.300 ;
      RECT 1478.830 0.700 1479.110 1511.300 ;
      RECT 1481.070 0.700 1481.350 1511.300 ;
      RECT 1483.310 0.700 1483.590 1511.300 ;
      RECT 1485.550 0.700 1485.830 1511.300 ;
      RECT 1487.790 0.700 1488.070 1511.300 ;
      RECT 1490.030 0.700 1490.310 1511.300 ;
      RECT 1492.270 0.700 1492.550 1511.300 ;
      RECT 1494.510 0.700 1494.790 1511.300 ;
      RECT 1496.750 0.700 1497.030 1511.300 ;
      RECT 1498.990 0.700 1499.270 1511.300 ;
      RECT 1501.230 0.700 1501.510 1511.300 ;
      RECT 1503.470 0.700 1503.750 1511.300 ;
      RECT 1505.710 0.700 1505.990 1511.300 ;
      RECT 1507.950 0.700 1508.230 1511.300 ;
      RECT 1510.190 0.700 1510.470 1511.300 ;
      RECT 1512.430 0.700 1512.710 1511.300 ;
      RECT 1514.670 0.700 1514.950 1511.300 ;
      RECT 1516.910 0.700 1517.190 1511.300 ;
      RECT 1519.150 0.700 1519.430 1511.300 ;
      RECT 1521.390 0.700 1521.670 1511.300 ;
      RECT 1523.630 0.700 1523.910 1511.300 ;
      RECT 1525.870 0.700 1526.150 1511.300 ;
      RECT 1528.110 0.700 1528.390 1511.300 ;
      RECT 1530.350 0.700 1530.630 1511.300 ;
      RECT 1532.590 0.700 1532.870 1511.300 ;
      RECT 1534.830 0.700 1535.110 1511.300 ;
      RECT 1537.070 0.700 1537.350 1511.300 ;
      RECT 1539.310 0.700 1539.590 1511.300 ;
      RECT 1541.550 0.700 1541.830 1511.300 ;
      RECT 1543.790 0.700 1544.070 1511.300 ;
      RECT 1546.030 0.700 1546.310 1511.300 ;
      RECT 1548.270 0.700 1548.550 1511.300 ;
      RECT 1550.510 0.700 1550.790 1511.300 ;
      RECT 1552.750 0.700 1553.030 1511.300 ;
      RECT 1554.990 0.700 1555.270 1511.300 ;
      RECT 1557.230 0.700 1557.510 1511.300 ;
      RECT 1559.470 0.700 1559.750 1511.300 ;
      RECT 1561.710 0.700 1561.990 1511.300 ;
      RECT 1563.950 0.700 1564.230 1511.300 ;
      RECT 1566.190 0.700 1566.470 1511.300 ;
      RECT 1568.430 0.700 1568.710 1511.300 ;
      RECT 1570.670 0.700 1570.950 1511.300 ;
      RECT 1572.910 0.700 1573.190 1511.300 ;
      RECT 1575.150 0.700 1575.430 1511.300 ;
      RECT 1577.390 0.700 1577.670 1511.300 ;
      RECT 1579.630 0.700 1579.910 1511.300 ;
      RECT 1581.870 0.700 1582.150 1511.300 ;
      RECT 1584.110 0.700 1584.390 1511.300 ;
      RECT 1586.350 0.700 1586.630 1511.300 ;
      RECT 1588.590 0.700 1588.870 1511.300 ;
      RECT 1590.830 0.700 1591.110 1511.300 ;
      RECT 1593.070 0.700 1593.350 1511.300 ;
      RECT 1595.310 0.700 1595.590 1511.300 ;
      RECT 1597.550 0.700 1597.830 1511.300 ;
      RECT 1599.790 0.700 1600.070 1511.300 ;
      RECT 1602.030 0.700 1602.310 1511.300 ;
      RECT 1604.270 0.700 1604.550 1511.300 ;
      RECT 1606.510 0.700 1606.790 1511.300 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 1609.300 1512.000 ;
    LAYER metal2 ;
    RECT 0 0 1609.300 1512.000 ;
    LAYER metal3 ;
    RECT 0 0 1609.300 1512.000 ;
    LAYER metal4 ;
    RECT 0 0 1609.300 1512.000 ;
    LAYER OVERLAP ;
    RECT 0 0 1609.300 1512.000 ;
  END
END fakeram_512x2048_1r1w

END LIBRARY
